module RecFNToIN( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@212294.2]
  input  [32:0] io_in, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@212295.4]
  input  [2:0]  io_roundingMode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@212295.4]
  input         io_signedOut, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@212295.4]
  output [31:0] io_out, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@212295.4]
  output [2:0]  io_intExceptionFlags // @[:freechips.rocketchip.system.DefaultRV32Config.fir@212295.4]
);
  wire  rawIn_isZero; // @[rawFloatFromRecFN.scala 51:54:freechips.rocketchip.system.DefaultRV32Config.fir@212300.4]
  wire  _T_4; // @[rawFloatFromRecFN.scala 52:54:freechips.rocketchip.system.DefaultRV32Config.fir@212302.4]
  wire  rawIn_isNaN; // @[rawFloatFromRecFN.scala 55:33:freechips.rocketchip.system.DefaultRV32Config.fir@212306.4]
  wire  _T_8; // @[rawFloatFromRecFN.scala 56:36:freechips.rocketchip.system.DefaultRV32Config.fir@212309.4]
  wire  rawIn_isInf; // @[rawFloatFromRecFN.scala 56:33:freechips.rocketchip.system.DefaultRV32Config.fir@212310.4]
  wire  rawIn_sign; // @[rawFloatFromRecFN.scala 58:25:freechips.rocketchip.system.DefaultRV32Config.fir@212313.4]
  wire [9:0] rawIn_sExp; // @[rawFloatFromRecFN.scala 59:27:freechips.rocketchip.system.DefaultRV32Config.fir@212315.4]
  wire  _T_12; // @[rawFloatFromRecFN.scala 60:39:freechips.rocketchip.system.DefaultRV32Config.fir@212317.4]
  wire [24:0] rawIn_sig; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@212320.4]
  wire  magGeOne; // @[RecFNToIN.scala 58:30:freechips.rocketchip.system.DefaultRV32Config.fir@212322.4]
  wire [7:0] posExp; // @[RecFNToIN.scala 59:28:freechips.rocketchip.system.DefaultRV32Config.fir@212323.4]
  wire  _T_16; // @[RecFNToIN.scala 60:27:freechips.rocketchip.system.DefaultRV32Config.fir@212324.4]
  wire  _T_17; // @[RecFNToIN.scala 60:47:freechips.rocketchip.system.DefaultRV32Config.fir@212325.4]
  wire  magJustBelowOne; // @[RecFNToIN.scala 60:37:freechips.rocketchip.system.DefaultRV32Config.fir@212326.4]
  wire  roundingMode_near_even; // @[RecFNToIN.scala 64:53:freechips.rocketchip.system.DefaultRV32Config.fir@212327.4]
  wire  roundingMode_min; // @[RecFNToIN.scala 66:53:freechips.rocketchip.system.DefaultRV32Config.fir@212329.4]
  wire  roundingMode_max; // @[RecFNToIN.scala 67:53:freechips.rocketchip.system.DefaultRV32Config.fir@212330.4]
  wire  roundingMode_near_maxMag; // @[RecFNToIN.scala 68:53:freechips.rocketchip.system.DefaultRV32Config.fir@212331.4]
  wire  roundingMode_odd; // @[RecFNToIN.scala 69:53:freechips.rocketchip.system.DefaultRV32Config.fir@212332.4]
  wire [23:0] _T_19; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@212334.4]
  wire [4:0] _T_21; // @[RecFNToIN.scala 81:16:freechips.rocketchip.system.DefaultRV32Config.fir@212336.4]
  wire [54:0] _GEN_0; // @[RecFNToIN.scala 80:50:freechips.rocketchip.system.DefaultRV32Config.fir@212337.4]
  wire [54:0] shiftedSig; // @[RecFNToIN.scala 80:50:freechips.rocketchip.system.DefaultRV32Config.fir@212337.4]
  wire  _T_24; // @[RecFNToIN.scala 86:69:freechips.rocketchip.system.DefaultRV32Config.fir@212340.4]
  wire [33:0] alignedSig; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@212341.4]
  wire [31:0] unroundedInt; // @[RecFNToIN.scala 87:54:freechips.rocketchip.system.DefaultRV32Config.fir@212342.4]
  wire  _T_27; // @[RecFNToIN.scala 89:57:freechips.rocketchip.system.DefaultRV32Config.fir@212345.4]
  wire  common_inexact; // @[RecFNToIN.scala 89:29:freechips.rocketchip.system.DefaultRV32Config.fir@212347.4]
  wire  _T_30; // @[RecFNToIN.scala 91:46:freechips.rocketchip.system.DefaultRV32Config.fir@212349.4]
  wire  _T_32; // @[RecFNToIN.scala 91:71:freechips.rocketchip.system.DefaultRV32Config.fir@212351.4]
  wire  _T_33; // @[RecFNToIN.scala 91:51:freechips.rocketchip.system.DefaultRV32Config.fir@212352.4]
  wire  _T_34; // @[RecFNToIN.scala 91:25:freechips.rocketchip.system.DefaultRV32Config.fir@212353.4]
  wire  _T_37; // @[RecFNToIN.scala 92:26:freechips.rocketchip.system.DefaultRV32Config.fir@212356.4]
  wire  roundIncr_near_even; // @[RecFNToIN.scala 91:78:freechips.rocketchip.system.DefaultRV32Config.fir@212357.4]
  wire  _T_39; // @[RecFNToIN.scala 93:43:freechips.rocketchip.system.DefaultRV32Config.fir@212359.4]
  wire  roundIncr_near_maxMag; // @[RecFNToIN.scala 93:61:freechips.rocketchip.system.DefaultRV32Config.fir@212360.4]
  wire  _T_40; // @[RecFNToIN.scala 95:35:freechips.rocketchip.system.DefaultRV32Config.fir@212361.4]
  wire  _T_41; // @[RecFNToIN.scala 96:35:freechips.rocketchip.system.DefaultRV32Config.fir@212362.4]
  wire  _T_42; // @[RecFNToIN.scala 95:61:freechips.rocketchip.system.DefaultRV32Config.fir@212363.4]
  wire  _T_43; // @[RecFNToIN.scala 97:28:freechips.rocketchip.system.DefaultRV32Config.fir@212364.4]
  wire  _T_44; // @[RecFNToIN.scala 98:26:freechips.rocketchip.system.DefaultRV32Config.fir@212365.4]
  wire  _T_45; // @[RecFNToIN.scala 97:49:freechips.rocketchip.system.DefaultRV32Config.fir@212366.4]
  wire  _T_46; // @[RecFNToIN.scala 96:61:freechips.rocketchip.system.DefaultRV32Config.fir@212367.4]
  wire  _T_47; // @[RecFNToIN.scala 99:31:freechips.rocketchip.system.DefaultRV32Config.fir@212368.4]
  wire  _T_48; // @[RecFNToIN.scala 99:43:freechips.rocketchip.system.DefaultRV32Config.fir@212369.4]
  wire  _T_49; // @[RecFNToIN.scala 99:27:freechips.rocketchip.system.DefaultRV32Config.fir@212370.4]
  wire  roundIncr; // @[RecFNToIN.scala 98:46:freechips.rocketchip.system.DefaultRV32Config.fir@212371.4]
  wire [31:0] _T_50; // @[RecFNToIN.scala 100:45:freechips.rocketchip.system.DefaultRV32Config.fir@212372.4]
  wire [31:0] complUnroundedInt; // @[RecFNToIN.scala 100:32:freechips.rocketchip.system.DefaultRV32Config.fir@212373.4]
  wire  _T_51; // @[RecFNToIN.scala 102:23:freechips.rocketchip.system.DefaultRV32Config.fir@212374.4]
  wire [31:0] _T_53; // @[RecFNToIN.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@212376.4]
  wire [31:0] _T_54; // @[RecFNToIN.scala 102:12:freechips.rocketchip.system.DefaultRV32Config.fir@212377.4]
  wire  _T_55; // @[RecFNToIN.scala 105:31:freechips.rocketchip.system.DefaultRV32Config.fir@212378.4]
  wire [31:0] _GEN_1; // @[RecFNToIN.scala 105:11:freechips.rocketchip.system.DefaultRV32Config.fir@212379.4]
  wire [31:0] roundedInt; // @[RecFNToIN.scala 105:11:freechips.rocketchip.system.DefaultRV32Config.fir@212379.4]
  wire  magGeOne_atOverflowEdge; // @[RecFNToIN.scala 107:43:freechips.rocketchip.system.DefaultRV32Config.fir@212380.4]
  wire  _T_57; // @[RecFNToIN.scala 110:56:freechips.rocketchip.system.DefaultRV32Config.fir@212382.4]
  wire  roundCarryBut2; // @[RecFNToIN.scala 110:61:freechips.rocketchip.system.DefaultRV32Config.fir@212383.4]
  wire  _T_58; // @[RecFNToIN.scala 113:21:freechips.rocketchip.system.DefaultRV32Config.fir@212384.4]
  wire  _T_60; // @[RecFNToIN.scala 117:60:freechips.rocketchip.system.DefaultRV32Config.fir@212386.4]
  wire  _T_61; // @[RecFNToIN.scala 117:64:freechips.rocketchip.system.DefaultRV32Config.fir@212387.4]
  wire  _T_62; // @[RecFNToIN.scala 116:49:freechips.rocketchip.system.DefaultRV32Config.fir@212388.4]
  wire  _T_63; // @[RecFNToIN.scala 119:38:freechips.rocketchip.system.DefaultRV32Config.fir@212389.4]
  wire  _T_64; // @[RecFNToIN.scala 119:62:freechips.rocketchip.system.DefaultRV32Config.fir@212390.4]
  wire  _T_65; // @[RecFNToIN.scala 118:49:freechips.rocketchip.system.DefaultRV32Config.fir@212391.4]
  wire  _T_66; // @[RecFNToIN.scala 115:24:freechips.rocketchip.system.DefaultRV32Config.fir@212392.4]
  wire  _T_68; // @[RecFNToIN.scala 122:50:freechips.rocketchip.system.DefaultRV32Config.fir@212394.4]
  wire  _T_69; // @[RecFNToIN.scala 123:57:freechips.rocketchip.system.DefaultRV32Config.fir@212395.4]
  wire  _T_70; // @[RecFNToIN.scala 121:32:freechips.rocketchip.system.DefaultRV32Config.fir@212396.4]
  wire  _T_71; // @[RecFNToIN.scala 114:20:freechips.rocketchip.system.DefaultRV32Config.fir@212397.4]
  wire  _T_72; // @[RecFNToIN.scala 113:40:freechips.rocketchip.system.DefaultRV32Config.fir@212398.4]
  wire  _T_73; // @[RecFNToIN.scala 125:13:freechips.rocketchip.system.DefaultRV32Config.fir@212399.4]
  wire  _T_74; // @[RecFNToIN.scala 125:27:freechips.rocketchip.system.DefaultRV32Config.fir@212400.4]
  wire  _T_75; // @[RecFNToIN.scala 125:41:freechips.rocketchip.system.DefaultRV32Config.fir@212401.4]
  wire  common_overflow; // @[RecFNToIN.scala 112:12:freechips.rocketchip.system.DefaultRV32Config.fir@212402.4]
  wire  invalidExc; // @[RecFNToIN.scala 130:34:freechips.rocketchip.system.DefaultRV32Config.fir@212403.4]
  wire  _T_76; // @[RecFNToIN.scala 131:20:freechips.rocketchip.system.DefaultRV32Config.fir@212404.4]
  wire  overflow; // @[RecFNToIN.scala 131:32:freechips.rocketchip.system.DefaultRV32Config.fir@212405.4]
  wire  _T_78; // @[RecFNToIN.scala 132:35:freechips.rocketchip.system.DefaultRV32Config.fir@212407.4]
  wire  _T_79; // @[RecFNToIN.scala 132:32:freechips.rocketchip.system.DefaultRV32Config.fir@212408.4]
  wire  inexact; // @[RecFNToIN.scala 132:52:freechips.rocketchip.system.DefaultRV32Config.fir@212409.4]
  wire  _T_80; // @[RecFNToIN.scala 134:19:freechips.rocketchip.system.DefaultRV32Config.fir@212410.4]
  wire  excSign; // @[RecFNToIN.scala 134:32:freechips.rocketchip.system.DefaultRV32Config.fir@212411.4]
  wire  _T_81; // @[RecFNToIN.scala 136:27:freechips.rocketchip.system.DefaultRV32Config.fir@212412.4]
  wire [31:0] _T_82; // @[RecFNToIN.scala 136:12:freechips.rocketchip.system.DefaultRV32Config.fir@212413.4]
  wire  _T_83; // @[RecFNToIN.scala 140:13:freechips.rocketchip.system.DefaultRV32Config.fir@212414.4]
  wire [30:0] _T_84; // @[RecFNToIN.scala 140:12:freechips.rocketchip.system.DefaultRV32Config.fir@212415.4]
  wire [31:0] _GEN_2; // @[RecFNToIN.scala 139:11:freechips.rocketchip.system.DefaultRV32Config.fir@212416.4]
  wire [31:0] excOut; // @[RecFNToIN.scala 139:11:freechips.rocketchip.system.DefaultRV32Config.fir@212416.4]
  wire  _T_85; // @[RecFNToIN.scala 142:30:freechips.rocketchip.system.DefaultRV32Config.fir@212417.4]
  wire [1:0] _T_87; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@212420.4]
  assign rawIn_isZero = io_in[31:29] == 3'h0; // @[rawFloatFromRecFN.scala 51:54:freechips.rocketchip.system.DefaultRV32Config.fir@212300.4]
  assign _T_4 = io_in[31:30] == 2'h3; // @[rawFloatFromRecFN.scala 52:54:freechips.rocketchip.system.DefaultRV32Config.fir@212302.4]
  assign rawIn_isNaN = _T_4 & io_in[29]; // @[rawFloatFromRecFN.scala 55:33:freechips.rocketchip.system.DefaultRV32Config.fir@212306.4]
  assign _T_8 = ~io_in[29]; // @[rawFloatFromRecFN.scala 56:36:freechips.rocketchip.system.DefaultRV32Config.fir@212309.4]
  assign rawIn_isInf = _T_4 & _T_8; // @[rawFloatFromRecFN.scala 56:33:freechips.rocketchip.system.DefaultRV32Config.fir@212310.4]
  assign rawIn_sign = io_in[32]; // @[rawFloatFromRecFN.scala 58:25:freechips.rocketchip.system.DefaultRV32Config.fir@212313.4]
  assign rawIn_sExp = {1'b0,$signed(io_in[31:23])}; // @[rawFloatFromRecFN.scala 59:27:freechips.rocketchip.system.DefaultRV32Config.fir@212315.4]
  assign _T_12 = ~rawIn_isZero; // @[rawFloatFromRecFN.scala 60:39:freechips.rocketchip.system.DefaultRV32Config.fir@212317.4]
  assign rawIn_sig = {1'h0,_T_12,io_in[22:0]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@212320.4]
  assign magGeOne = rawIn_sExp[8]; // @[RecFNToIN.scala 58:30:freechips.rocketchip.system.DefaultRV32Config.fir@212322.4]
  assign posExp = rawIn_sExp[7:0]; // @[RecFNToIN.scala 59:28:freechips.rocketchip.system.DefaultRV32Config.fir@212323.4]
  assign _T_16 = ~magGeOne; // @[RecFNToIN.scala 60:27:freechips.rocketchip.system.DefaultRV32Config.fir@212324.4]
  assign _T_17 = &posExp; // @[RecFNToIN.scala 60:47:freechips.rocketchip.system.DefaultRV32Config.fir@212325.4]
  assign magJustBelowOne = _T_16 & _T_17; // @[RecFNToIN.scala 60:37:freechips.rocketchip.system.DefaultRV32Config.fir@212326.4]
  assign roundingMode_near_even = io_roundingMode == 3'h0; // @[RecFNToIN.scala 64:53:freechips.rocketchip.system.DefaultRV32Config.fir@212327.4]
  assign roundingMode_min = io_roundingMode == 3'h2; // @[RecFNToIN.scala 66:53:freechips.rocketchip.system.DefaultRV32Config.fir@212329.4]
  assign roundingMode_max = io_roundingMode == 3'h3; // @[RecFNToIN.scala 67:53:freechips.rocketchip.system.DefaultRV32Config.fir@212330.4]
  assign roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RecFNToIN.scala 68:53:freechips.rocketchip.system.DefaultRV32Config.fir@212331.4]
  assign roundingMode_odd = io_roundingMode == 3'h6; // @[RecFNToIN.scala 69:53:freechips.rocketchip.system.DefaultRV32Config.fir@212332.4]
  assign _T_19 = {magGeOne,rawIn_sig[22:0]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@212334.4]
  assign _T_21 = magGeOne ? rawIn_sExp[4:0] : 5'h0; // @[RecFNToIN.scala 81:16:freechips.rocketchip.system.DefaultRV32Config.fir@212336.4]
  assign _GEN_0 = {{31'd0}, _T_19}; // @[RecFNToIN.scala 80:50:freechips.rocketchip.system.DefaultRV32Config.fir@212337.4]
  assign shiftedSig = _GEN_0 << _T_21; // @[RecFNToIN.scala 80:50:freechips.rocketchip.system.DefaultRV32Config.fir@212337.4]
  assign _T_24 = |shiftedSig[21:0]; // @[RecFNToIN.scala 86:69:freechips.rocketchip.system.DefaultRV32Config.fir@212340.4]
  assign alignedSig = {shiftedSig[54:22],_T_24}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@212341.4]
  assign unroundedInt = alignedSig[33:2]; // @[RecFNToIN.scala 87:54:freechips.rocketchip.system.DefaultRV32Config.fir@212342.4]
  assign _T_27 = |alignedSig[1:0]; // @[RecFNToIN.scala 89:57:freechips.rocketchip.system.DefaultRV32Config.fir@212345.4]
  assign common_inexact = magGeOne ? _T_27 : _T_12; // @[RecFNToIN.scala 89:29:freechips.rocketchip.system.DefaultRV32Config.fir@212347.4]
  assign _T_30 = &alignedSig[2:1]; // @[RecFNToIN.scala 91:46:freechips.rocketchip.system.DefaultRV32Config.fir@212349.4]
  assign _T_32 = &alignedSig[1:0]; // @[RecFNToIN.scala 91:71:freechips.rocketchip.system.DefaultRV32Config.fir@212351.4]
  assign _T_33 = _T_30 | _T_32; // @[RecFNToIN.scala 91:51:freechips.rocketchip.system.DefaultRV32Config.fir@212352.4]
  assign _T_34 = magGeOne & _T_33; // @[RecFNToIN.scala 91:25:freechips.rocketchip.system.DefaultRV32Config.fir@212353.4]
  assign _T_37 = magJustBelowOne & _T_27; // @[RecFNToIN.scala 92:26:freechips.rocketchip.system.DefaultRV32Config.fir@212356.4]
  assign roundIncr_near_even = _T_34 | _T_37; // @[RecFNToIN.scala 91:78:freechips.rocketchip.system.DefaultRV32Config.fir@212357.4]
  assign _T_39 = magGeOne & alignedSig[1]; // @[RecFNToIN.scala 93:43:freechips.rocketchip.system.DefaultRV32Config.fir@212359.4]
  assign roundIncr_near_maxMag = _T_39 | magJustBelowOne; // @[RecFNToIN.scala 93:61:freechips.rocketchip.system.DefaultRV32Config.fir@212360.4]
  assign _T_40 = roundingMode_near_even & roundIncr_near_even; // @[RecFNToIN.scala 95:35:freechips.rocketchip.system.DefaultRV32Config.fir@212361.4]
  assign _T_41 = roundingMode_near_maxMag & roundIncr_near_maxMag; // @[RecFNToIN.scala 96:35:freechips.rocketchip.system.DefaultRV32Config.fir@212362.4]
  assign _T_42 = _T_40 | _T_41; // @[RecFNToIN.scala 95:61:freechips.rocketchip.system.DefaultRV32Config.fir@212363.4]
  assign _T_43 = roundingMode_min | roundingMode_odd; // @[RecFNToIN.scala 97:28:freechips.rocketchip.system.DefaultRV32Config.fir@212364.4]
  assign _T_44 = rawIn_sign & common_inexact; // @[RecFNToIN.scala 98:26:freechips.rocketchip.system.DefaultRV32Config.fir@212365.4]
  assign _T_45 = _T_43 & _T_44; // @[RecFNToIN.scala 97:49:freechips.rocketchip.system.DefaultRV32Config.fir@212366.4]
  assign _T_46 = _T_42 | _T_45; // @[RecFNToIN.scala 96:61:freechips.rocketchip.system.DefaultRV32Config.fir@212367.4]
  assign _T_47 = ~rawIn_sign; // @[RecFNToIN.scala 99:31:freechips.rocketchip.system.DefaultRV32Config.fir@212368.4]
  assign _T_48 = _T_47 & common_inexact; // @[RecFNToIN.scala 99:43:freechips.rocketchip.system.DefaultRV32Config.fir@212369.4]
  assign _T_49 = roundingMode_max & _T_48; // @[RecFNToIN.scala 99:27:freechips.rocketchip.system.DefaultRV32Config.fir@212370.4]
  assign roundIncr = _T_46 | _T_49; // @[RecFNToIN.scala 98:46:freechips.rocketchip.system.DefaultRV32Config.fir@212371.4]
  assign _T_50 = ~unroundedInt; // @[RecFNToIN.scala 100:45:freechips.rocketchip.system.DefaultRV32Config.fir@212372.4]
  assign complUnroundedInt = rawIn_sign ? _T_50 : unroundedInt; // @[RecFNToIN.scala 100:32:freechips.rocketchip.system.DefaultRV32Config.fir@212373.4]
  assign _T_51 = roundIncr ^ rawIn_sign; // @[RecFNToIN.scala 102:23:freechips.rocketchip.system.DefaultRV32Config.fir@212374.4]
  assign _T_53 = complUnroundedInt + 32'h1; // @[RecFNToIN.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@212376.4]
  assign _T_54 = _T_51 ? _T_53 : complUnroundedInt; // @[RecFNToIN.scala 102:12:freechips.rocketchip.system.DefaultRV32Config.fir@212377.4]
  assign _T_55 = roundingMode_odd & common_inexact; // @[RecFNToIN.scala 105:31:freechips.rocketchip.system.DefaultRV32Config.fir@212378.4]
  assign _GEN_1 = {{31'd0}, _T_55}; // @[RecFNToIN.scala 105:11:freechips.rocketchip.system.DefaultRV32Config.fir@212379.4]
  assign roundedInt = _T_54 | _GEN_1; // @[RecFNToIN.scala 105:11:freechips.rocketchip.system.DefaultRV32Config.fir@212379.4]
  assign magGeOne_atOverflowEdge = posExp == 8'h1f; // @[RecFNToIN.scala 107:43:freechips.rocketchip.system.DefaultRV32Config.fir@212380.4]
  assign _T_57 = &unroundedInt[29:0]; // @[RecFNToIN.scala 110:56:freechips.rocketchip.system.DefaultRV32Config.fir@212382.4]
  assign roundCarryBut2 = _T_57 & roundIncr; // @[RecFNToIN.scala 110:61:freechips.rocketchip.system.DefaultRV32Config.fir@212383.4]
  assign _T_58 = posExp >= 8'h20; // @[RecFNToIN.scala 113:21:freechips.rocketchip.system.DefaultRV32Config.fir@212384.4]
  assign _T_60 = |unroundedInt[30:0]; // @[RecFNToIN.scala 117:60:freechips.rocketchip.system.DefaultRV32Config.fir@212386.4]
  assign _T_61 = _T_60 | roundIncr; // @[RecFNToIN.scala 117:64:freechips.rocketchip.system.DefaultRV32Config.fir@212387.4]
  assign _T_62 = magGeOne_atOverflowEdge & _T_61; // @[RecFNToIN.scala 116:49:freechips.rocketchip.system.DefaultRV32Config.fir@212388.4]
  assign _T_63 = posExp == 8'h1e; // @[RecFNToIN.scala 119:38:freechips.rocketchip.system.DefaultRV32Config.fir@212389.4]
  assign _T_64 = _T_63 & roundCarryBut2; // @[RecFNToIN.scala 119:62:freechips.rocketchip.system.DefaultRV32Config.fir@212390.4]
  assign _T_65 = magGeOne_atOverflowEdge | _T_64; // @[RecFNToIN.scala 118:49:freechips.rocketchip.system.DefaultRV32Config.fir@212391.4]
  assign _T_66 = rawIn_sign ? _T_62 : _T_65; // @[RecFNToIN.scala 115:24:freechips.rocketchip.system.DefaultRV32Config.fir@212392.4]
  assign _T_68 = magGeOne_atOverflowEdge & unroundedInt[30]; // @[RecFNToIN.scala 122:50:freechips.rocketchip.system.DefaultRV32Config.fir@212394.4]
  assign _T_69 = _T_68 & roundCarryBut2; // @[RecFNToIN.scala 123:57:freechips.rocketchip.system.DefaultRV32Config.fir@212395.4]
  assign _T_70 = rawIn_sign | _T_69; // @[RecFNToIN.scala 121:32:freechips.rocketchip.system.DefaultRV32Config.fir@212396.4]
  assign _T_71 = io_signedOut ? _T_66 : _T_70; // @[RecFNToIN.scala 114:20:freechips.rocketchip.system.DefaultRV32Config.fir@212397.4]
  assign _T_72 = _T_58 | _T_71; // @[RecFNToIN.scala 113:40:freechips.rocketchip.system.DefaultRV32Config.fir@212398.4]
  assign _T_73 = ~io_signedOut; // @[RecFNToIN.scala 125:13:freechips.rocketchip.system.DefaultRV32Config.fir@212399.4]
  assign _T_74 = _T_73 & rawIn_sign; // @[RecFNToIN.scala 125:27:freechips.rocketchip.system.DefaultRV32Config.fir@212400.4]
  assign _T_75 = _T_74 & roundIncr; // @[RecFNToIN.scala 125:41:freechips.rocketchip.system.DefaultRV32Config.fir@212401.4]
  assign common_overflow = magGeOne ? _T_72 : _T_75; // @[RecFNToIN.scala 112:12:freechips.rocketchip.system.DefaultRV32Config.fir@212402.4]
  assign invalidExc = rawIn_isNaN | rawIn_isInf; // @[RecFNToIN.scala 130:34:freechips.rocketchip.system.DefaultRV32Config.fir@212403.4]
  assign _T_76 = ~invalidExc; // @[RecFNToIN.scala 131:20:freechips.rocketchip.system.DefaultRV32Config.fir@212404.4]
  assign overflow = _T_76 & common_overflow; // @[RecFNToIN.scala 131:32:freechips.rocketchip.system.DefaultRV32Config.fir@212405.4]
  assign _T_78 = ~common_overflow; // @[RecFNToIN.scala 132:35:freechips.rocketchip.system.DefaultRV32Config.fir@212407.4]
  assign _T_79 = _T_76 & _T_78; // @[RecFNToIN.scala 132:32:freechips.rocketchip.system.DefaultRV32Config.fir@212408.4]
  assign inexact = _T_79 & common_inexact; // @[RecFNToIN.scala 132:52:freechips.rocketchip.system.DefaultRV32Config.fir@212409.4]
  assign _T_80 = ~rawIn_isNaN; // @[RecFNToIN.scala 134:19:freechips.rocketchip.system.DefaultRV32Config.fir@212410.4]
  assign excSign = _T_80 & rawIn_sign; // @[RecFNToIN.scala 134:32:freechips.rocketchip.system.DefaultRV32Config.fir@212411.4]
  assign _T_81 = io_signedOut == excSign; // @[RecFNToIN.scala 136:27:freechips.rocketchip.system.DefaultRV32Config.fir@212412.4]
  assign _T_82 = _T_81 ? 32'h80000000 : 32'h0; // @[RecFNToIN.scala 136:12:freechips.rocketchip.system.DefaultRV32Config.fir@212413.4]
  assign _T_83 = ~excSign; // @[RecFNToIN.scala 140:13:freechips.rocketchip.system.DefaultRV32Config.fir@212414.4]
  assign _T_84 = _T_83 ? 31'h7fffffff : 31'h0; // @[RecFNToIN.scala 140:12:freechips.rocketchip.system.DefaultRV32Config.fir@212415.4]
  assign _GEN_2 = {{1'd0}, _T_84}; // @[RecFNToIN.scala 139:11:freechips.rocketchip.system.DefaultRV32Config.fir@212416.4]
  assign excOut = _T_82 | _GEN_2; // @[RecFNToIN.scala 139:11:freechips.rocketchip.system.DefaultRV32Config.fir@212416.4]
  assign _T_85 = invalidExc | common_overflow; // @[RecFNToIN.scala 142:30:freechips.rocketchip.system.DefaultRV32Config.fir@212417.4]
  assign _T_87 = {invalidExc,overflow}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@212420.4]
  assign io_out = _T_85 ? excOut : roundedInt; // @[RecFNToIN.scala 142:12:freechips.rocketchip.system.DefaultRV32Config.fir@212419.4]
  assign io_intExceptionFlags = {_T_87,inexact}; // @[RecFNToIN.scala 143:26:freechips.rocketchip.system.DefaultRV32Config.fir@212422.4]
endmodule
