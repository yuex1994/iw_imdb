module OptimizationBarrier_117( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214465.2]
  input  [2:0] io_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214468.4]
  output [2:0] io_y // @[:freechips.rocketchip.system.DefaultRV32Config.fir@214468.4]
);
  assign io_y = io_x; // @[package.scala 236:12:freechips.rocketchip.system.DefaultRV32Config.fir@214473.4]
endmodule
