module RVCExpander( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@215557.2]
  input  [31:0] io_in, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@215560.4]
  output [31:0] io_out_bits, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@215560.4]
  output [4:0]  io_out_rd, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@215560.4]
  output [4:0]  io_out_rs1, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@215560.4]
  output [4:0]  io_out_rs2, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@215560.4]
  output [4:0]  io_out_rs3, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@215560.4]
  output        io_rvc // @[:freechips.rocketchip.system.DefaultRV32Config.fir@215560.4]
);
  wire  _T_3; // @[RVC.scala 54:29:freechips.rocketchip.system.DefaultRV32Config.fir@215566.4]
  wire [6:0] _T_4; // @[RVC.scala 54:20:freechips.rocketchip.system.DefaultRV32Config.fir@215567.4]
  wire [4:0] _T_14; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215577.4]
  wire [29:0] _T_18; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215581.4]
  wire [7:0] _T_28; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215596.4]
  wire [4:0] _T_30; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215598.4]
  wire [27:0] _T_36; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215604.4]
  wire [6:0] _T_50; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215623.4]
  wire [26:0] _T_58; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215631.4]
  wire [26:0] _T_80; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215658.4]
  wire [26:0] _T_111; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215694.4]
  wire [27:0] _T_138; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215726.4]
  wire [26:0] _T_169; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215762.4]
  wire [26:0] _T_200; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215798.4]
  wire [6:0] _T_211; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@215814.4]
  wire [11:0] _T_213; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215816.4]
  wire [31:0] _T_219; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215822.4]
  wire [9:0] _T_228; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@215836.4]
  wire [20:0] _T_243; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215851.4]
  wire [31:0] _T_306; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215914.4]
  wire [31:0] _T_321; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215934.4]
  wire  _T_332; // @[RVC.scala 91:29:freechips.rocketchip.system.DefaultRV32Config.fir@215950.4]
  wire [6:0] _T_333; // @[RVC.scala 91:20:freechips.rocketchip.system.DefaultRV32Config.fir@215951.4]
  wire [14:0] _T_336; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@215954.4]
  wire [31:0] _T_339; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215957.4]
  wire [31:0] _T_343; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215961.4]
  wire  _T_351; // @[RVC.scala 93:14:freechips.rocketchip.system.DefaultRV32Config.fir@215974.4]
  wire  _T_353; // @[RVC.scala 93:27:freechips.rocketchip.system.DefaultRV32Config.fir@215976.4]
  wire  _T_354; // @[RVC.scala 93:21:freechips.rocketchip.system.DefaultRV32Config.fir@215977.4]
  wire [6:0] _T_361; // @[RVC.scala 87:20:freechips.rocketchip.system.DefaultRV32Config.fir@215984.4]
  wire [2:0] _T_364; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@215987.4]
  wire [31:0] _T_379; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216002.4]
  wire [31:0] _T_386_bits; // @[RVC.scala 93:10:freechips.rocketchip.system.DefaultRV32Config.fir@216014.4]
  wire [4:0] _T_386_rd; // @[RVC.scala 93:10:freechips.rocketchip.system.DefaultRV32Config.fir@216014.4]
  wire [4:0] _T_386_rs2; // @[RVC.scala 93:10:freechips.rocketchip.system.DefaultRV32Config.fir@216014.4]
  wire [4:0] _T_386_rs3; // @[RVC.scala 93:10:freechips.rocketchip.system.DefaultRV32Config.fir@216014.4]
  wire [25:0] _T_397; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216025.4]
  wire [30:0] _GEN_0; // @[RVC.scala 100:23:freechips.rocketchip.system.DefaultRV32Config.fir@216037.4]
  wire [30:0] _T_409; // @[RVC.scala 100:23:freechips.rocketchip.system.DefaultRV32Config.fir@216037.4]
  wire [31:0] _T_422; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216050.4]
  wire [2:0] _T_425; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216053.4]
  wire  _T_426; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216054.4]
  wire [2:0] _T_427; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216055.4]
  wire  _T_428; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216056.4]
  wire [2:0] _T_429; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216057.4]
  wire  _T_430; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216058.4]
  wire [2:0] _T_431; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216059.4]
  wire  _T_432; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216060.4]
  wire [2:0] _T_433; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216061.4]
  wire  _T_434; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216062.4]
  wire [2:0] _T_435; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216063.4]
  wire  _T_436; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216064.4]
  wire [2:0] _T_437; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216065.4]
  wire  _T_438; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216066.4]
  wire [2:0] _T_439; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216067.4]
  wire  _T_441; // @[RVC.scala 104:30:freechips.rocketchip.system.DefaultRV32Config.fir@216069.4]
  wire [30:0] _T_442; // @[RVC.scala 104:22:freechips.rocketchip.system.DefaultRV32Config.fir@216070.4]
  wire [6:0] _T_444; // @[RVC.scala 105:22:freechips.rocketchip.system.DefaultRV32Config.fir@216072.4]
  wire [24:0] _T_454; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216082.4]
  wire [30:0] _GEN_1; // @[RVC.scala 106:43:freechips.rocketchip.system.DefaultRV32Config.fir@216083.4]
  wire [30:0] _T_455; // @[RVC.scala 106:43:freechips.rocketchip.system.DefaultRV32Config.fir@216083.4]
  wire  _T_457; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216085.4]
  wire [30:0] _T_458; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216086.4]
  wire  _T_459; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216087.4]
  wire [31:0] _T_460; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216088.4]
  wire  _T_461; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216089.4]
  wire [31:0] _T_462; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216090.4]
  wire [31:0] _T_551; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216184.4]
  wire [4:0] _T_560; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@216198.4]
  wire [12:0] _T_569; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216207.4]
  wire [31:0] _T_618; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216256.4]
  wire [31:0] _T_685; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216328.4]
  wire  _T_691; // @[RVC.scala 114:27:freechips.rocketchip.system.DefaultRV32Config.fir@216339.4]
  wire [6:0] _T_692; // @[RVC.scala 114:23:freechips.rocketchip.system.DefaultRV32Config.fir@216340.4]
  wire [25:0] _T_701; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216349.4]
  wire [28:0] _T_717; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216370.4]
  wire [27:0] _T_732; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216390.4]
  wire [27:0] _T_747; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216410.4]
  wire [24:0] _T_757; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216425.4]
  wire [24:0] _T_768; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216441.4]
  wire [24:0] _T_779; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216457.4]
  wire [24:0] _T_781; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216459.4]
  wire [24:0] _T_784; // @[RVC.scala 135:33:freechips.rocketchip.system.DefaultRV32Config.fir@216462.4]
  wire  _T_790; // @[RVC.scala 136:27:freechips.rocketchip.system.DefaultRV32Config.fir@216473.4]
  wire [31:0] _T_761_bits; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@216429.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@216430.4]
  wire [31:0] _T_788_bits; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@216466.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@216467.4]
  wire [31:0] _T_791_bits; // @[RVC.scala 136:22:freechips.rocketchip.system.DefaultRV32Config.fir@216474.4]
  wire [4:0] _T_791_rd; // @[RVC.scala 136:22:freechips.rocketchip.system.DefaultRV32Config.fir@216474.4]
  wire [4:0] _T_791_rs1; // @[RVC.scala 136:22:freechips.rocketchip.system.DefaultRV32Config.fir@216474.4]
  wire [4:0] _T_791_rs2; // @[RVC.scala 136:22:freechips.rocketchip.system.DefaultRV32Config.fir@216474.4]
  wire [4:0] _T_791_rs3; // @[RVC.scala 136:22:freechips.rocketchip.system.DefaultRV32Config.fir@216474.4]
  wire [24:0] _T_797; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216480.4]
  wire [24:0] _T_799; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216482.4]
  wire [24:0] _T_800; // @[RVC.scala 138:46:freechips.rocketchip.system.DefaultRV32Config.fir@216483.4]
  wire [24:0] _T_803; // @[RVC.scala 139:33:freechips.rocketchip.system.DefaultRV32Config.fir@216486.4]
  wire [31:0] _T_773_bits; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@216446.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@216447.4]
  wire [31:0] _T_807_bits; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@216490.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@216491.4]
  wire [31:0] _T_810_bits; // @[RVC.scala 140:25:freechips.rocketchip.system.DefaultRV32Config.fir@216498.4]
  wire [4:0] _T_810_rd; // @[RVC.scala 140:25:freechips.rocketchip.system.DefaultRV32Config.fir@216498.4]
  wire [4:0] _T_810_rs1; // @[RVC.scala 140:25:freechips.rocketchip.system.DefaultRV32Config.fir@216498.4]
  wire [31:0] _T_812_bits; // @[RVC.scala 141:10:freechips.rocketchip.system.DefaultRV32Config.fir@216500.4]
  wire [4:0] _T_812_rd; // @[RVC.scala 141:10:freechips.rocketchip.system.DefaultRV32Config.fir@216500.4]
  wire [4:0] _T_812_rs1; // @[RVC.scala 141:10:freechips.rocketchip.system.DefaultRV32Config.fir@216500.4]
  wire [4:0] _T_812_rs2; // @[RVC.scala 141:10:freechips.rocketchip.system.DefaultRV32Config.fir@216500.4]
  wire [4:0] _T_812_rs3; // @[RVC.scala 141:10:freechips.rocketchip.system.DefaultRV32Config.fir@216500.4]
  wire [8:0] _T_816; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216504.4]
  wire [28:0] _T_828; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216516.4]
  wire [7:0] _T_836; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216529.4]
  wire [27:0] _T_848; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216541.4]
  wire [27:0] _T_868; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216566.4]
  wire [4:0] _T_915; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216658.4]
  wire  _T_916; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216659.4]
  wire [31:0] _T_44_bits; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@215612.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@215613.4]
  wire [31:0] _T_24_bits; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@215587.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@215588.4]
  wire [31:0] _T_917_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216660.4]
  wire [4:0] _T_917_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216660.4]
  wire [4:0] _T_917_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216660.4]
  wire [4:0] _T_917_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216660.4]
  wire  _T_918; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216661.4]
  wire [31:0] _T_66_bits; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@215639.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@215640.4]
  wire [31:0] _T_919_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216662.4]
  wire [4:0] _T_919_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216662.4]
  wire [4:0] _T_919_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216662.4]
  wire [4:0] _T_919_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216662.4]
  wire  _T_920; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216663.4]
  wire [31:0] _T_88_bits; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@215666.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@215667.4]
  wire [31:0] _T_921_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216664.4]
  wire [4:0] _T_921_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216664.4]
  wire [4:0] _T_921_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216664.4]
  wire [4:0] _T_921_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216664.4]
  wire  _T_922; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216665.4]
  wire [31:0] _T_119_bits; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@215702.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@215703.4]
  wire [31:0] _T_923_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216666.4]
  wire [4:0] _T_923_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216666.4]
  wire [4:0] _T_923_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216666.4]
  wire [4:0] _T_923_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216666.4]
  wire  _T_924; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216667.4]
  wire [31:0] _T_146_bits; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@215734.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@215735.4]
  wire [31:0] _T_925_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216668.4]
  wire [4:0] _T_925_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216668.4]
  wire [4:0] _T_925_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216668.4]
  wire [4:0] _T_925_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216668.4]
  wire  _T_926; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216669.4]
  wire [31:0] _T_177_bits; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@215770.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@215771.4]
  wire [31:0] _T_927_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216670.4]
  wire [4:0] _T_927_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216670.4]
  wire [4:0] _T_927_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216670.4]
  wire [4:0] _T_927_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216670.4]
  wire  _T_928; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216671.4]
  wire [31:0] _T_208_bits; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@215806.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@215807.4]
  wire [31:0] _T_929_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216672.4]
  wire [4:0] _T_929_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216672.4]
  wire [4:0] _T_929_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216672.4]
  wire [4:0] _T_929_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216672.4]
  wire  _T_930; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216673.4]
  wire [31:0] _T_931_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216674.4]
  wire [4:0] _T_931_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216674.4]
  wire [4:0] _T_931_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216674.4]
  wire [4:0] _T_931_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216674.4]
  wire [4:0] _T_931_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216674.4]
  wire  _T_932; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216675.4]
  wire [31:0] _T_933_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216676.4]
  wire [4:0] _T_933_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216676.4]
  wire [4:0] _T_933_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216676.4]
  wire [4:0] _T_933_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216676.4]
  wire [4:0] _T_933_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216676.4]
  wire  _T_934; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216677.4]
  wire [31:0] _T_935_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216678.4]
  wire [4:0] _T_935_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216678.4]
  wire [4:0] _T_935_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216678.4]
  wire [4:0] _T_935_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216678.4]
  wire [4:0] _T_935_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216678.4]
  wire  _T_936; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216679.4]
  wire [31:0] _T_937_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216680.4]
  wire [4:0] _T_937_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216680.4]
  wire [4:0] _T_937_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216680.4]
  wire [4:0] _T_937_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216680.4]
  wire [4:0] _T_937_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216680.4]
  wire  _T_938; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216681.4]
  wire [31:0] _T_939_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216682.4]
  wire [4:0] _T_939_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216682.4]
  wire [4:0] _T_939_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216682.4]
  wire [4:0] _T_939_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216682.4]
  wire [4:0] _T_939_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216682.4]
  wire  _T_940; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216683.4]
  wire [31:0] _T_941_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216684.4]
  wire [4:0] _T_941_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216684.4]
  wire [4:0] _T_941_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216684.4]
  wire [4:0] _T_941_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216684.4]
  wire [4:0] _T_941_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216684.4]
  wire  _T_942; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216685.4]
  wire [31:0] _T_943_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216686.4]
  wire [4:0] _T_943_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216686.4]
  wire [4:0] _T_943_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216686.4]
  wire [4:0] _T_943_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216686.4]
  wire [4:0] _T_943_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216686.4]
  wire  _T_944; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216687.4]
  wire [31:0] _T_945_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216688.4]
  wire [4:0] _T_945_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216688.4]
  wire [4:0] _T_945_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216688.4]
  wire [4:0] _T_945_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216688.4]
  wire [4:0] _T_945_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216688.4]
  wire  _T_946; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216689.4]
  wire [31:0] _T_706_bits; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@216354.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@216355.4]
  wire [31:0] _T_947_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216690.4]
  wire [4:0] _T_947_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216690.4]
  wire [4:0] _T_947_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216690.4]
  wire [4:0] _T_947_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216690.4]
  wire [4:0] _T_947_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216690.4]
  wire  _T_948; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216691.4]
  wire [31:0] _T_721_bits; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@216374.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@216375.4]
  wire [31:0] _T_949_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216692.4]
  wire [4:0] _T_949_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216692.4]
  wire [4:0] _T_949_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216692.4]
  wire [4:0] _T_949_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216692.4]
  wire [4:0] _T_949_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216692.4]
  wire  _T_950; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216693.4]
  wire [31:0] _T_736_bits; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@216394.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@216395.4]
  wire [31:0] _T_951_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216694.4]
  wire [4:0] _T_951_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216694.4]
  wire [4:0] _T_951_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216694.4]
  wire [4:0] _T_951_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216694.4]
  wire [4:0] _T_951_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216694.4]
  wire  _T_952; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216695.4]
  wire [31:0] _T_751_bits; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@216414.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@216415.4]
  wire [31:0] _T_953_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216696.4]
  wire [4:0] _T_953_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216696.4]
  wire [4:0] _T_953_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216696.4]
  wire [4:0] _T_953_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216696.4]
  wire [4:0] _T_953_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216696.4]
  wire  _T_954; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216697.4]
  wire [31:0] _T_955_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216698.4]
  wire [4:0] _T_955_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216698.4]
  wire [4:0] _T_955_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216698.4]
  wire [4:0] _T_955_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216698.4]
  wire [4:0] _T_955_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216698.4]
  wire  _T_956; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216699.4]
  wire [31:0] _T_832_bits; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@216520.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@216521.4]
  wire [31:0] _T_957_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216700.4]
  wire [4:0] _T_957_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216700.4]
  wire [4:0] _T_957_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216700.4]
  wire [4:0] _T_957_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216700.4]
  wire [4:0] _T_957_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216700.4]
  wire  _T_958; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216701.4]
  wire [31:0] _T_852_bits; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@216545.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@216546.4]
  wire [31:0] _T_959_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216702.4]
  wire [4:0] _T_959_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216702.4]
  wire [4:0] _T_959_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216702.4]
  wire [4:0] _T_959_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216702.4]
  wire [4:0] _T_959_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216702.4]
  wire  _T_960; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216703.4]
  wire [31:0] _T_872_bits; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@216570.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@216571.4]
  wire [31:0] _T_961_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216704.4]
  wire [4:0] _T_961_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216704.4]
  wire [4:0] _T_961_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216704.4]
  wire [4:0] _T_961_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216704.4]
  wire [4:0] _T_961_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216704.4]
  wire  _T_962; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216705.4]
  wire [31:0] _T_963_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216706.4]
  wire [4:0] _T_963_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216706.4]
  wire [4:0] _T_963_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216706.4]
  wire [4:0] _T_963_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216706.4]
  wire [4:0] _T_963_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216706.4]
  wire  _T_964; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216707.4]
  wire [31:0] _T_965_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216708.4]
  wire [4:0] _T_965_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216708.4]
  wire [4:0] _T_965_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216708.4]
  wire [4:0] _T_965_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216708.4]
  wire [4:0] _T_965_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216708.4]
  wire  _T_966; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216709.4]
  wire [31:0] _T_967_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216710.4]
  wire [4:0] _T_967_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216710.4]
  wire [4:0] _T_967_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216710.4]
  wire [4:0] _T_967_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216710.4]
  wire [4:0] _T_967_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216710.4]
  wire  _T_968; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216711.4]
  wire [31:0] _T_969_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216712.4]
  wire [4:0] _T_969_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216712.4]
  wire [4:0] _T_969_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216712.4]
  wire [4:0] _T_969_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216712.4]
  wire [4:0] _T_969_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216712.4]
  wire  _T_970; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216713.4]
  wire [31:0] _T_971_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216714.4]
  wire [4:0] _T_971_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216714.4]
  wire [4:0] _T_971_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216714.4]
  wire [4:0] _T_971_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216714.4]
  wire [4:0] _T_971_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216714.4]
  wire  _T_972; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216715.4]
  wire [31:0] _T_973_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216716.4]
  wire [4:0] _T_973_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216716.4]
  wire [4:0] _T_973_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216716.4]
  wire [4:0] _T_973_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216716.4]
  wire [4:0] _T_973_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216716.4]
  wire  _T_974; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216717.4]
  wire [31:0] _T_975_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216718.4]
  wire [4:0] _T_975_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216718.4]
  wire [4:0] _T_975_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216718.4]
  wire [4:0] _T_975_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216718.4]
  wire [4:0] _T_975_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216718.4]
  wire  _T_976; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216719.4]
  assign _T_3 = |io_in[12:5]; // @[RVC.scala 54:29:freechips.rocketchip.system.DefaultRV32Config.fir@215566.4]
  assign _T_4 = _T_3 ? 7'h13 : 7'h1f; // @[RVC.scala 54:20:freechips.rocketchip.system.DefaultRV32Config.fir@215567.4]
  assign _T_14 = {2'h1,io_in[4:2]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215577.4]
  assign _T_18 = {io_in[10:7],io_in[12:11],io_in[5],io_in[6],2'h0,5'h2,3'h0,2'h1,io_in[4:2],_T_4}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215581.4]
  assign _T_28 = {io_in[6:5],io_in[12:10],3'h0}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215596.4]
  assign _T_30 = {2'h1,io_in[9:7]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215598.4]
  assign _T_36 = {io_in[6:5],io_in[12:10],3'h0,2'h1,io_in[9:7],3'h3,2'h1,io_in[4:2],7'h7}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215604.4]
  assign _T_50 = {io_in[5],io_in[12:10],io_in[6],2'h0}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215623.4]
  assign _T_58 = {io_in[5],io_in[12:10],io_in[6],2'h0,2'h1,io_in[9:7],3'h2,2'h1,io_in[4:2],7'h3}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215631.4]
  assign _T_80 = {io_in[5],io_in[12:10],io_in[6],2'h0,2'h1,io_in[9:7],3'h2,2'h1,io_in[4:2],7'h7}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215658.4]
  assign _T_111 = {_T_50[6:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h2,_T_50[4:0],7'h3f}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215694.4]
  assign _T_138 = {_T_28[7:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h3,_T_28[4:0],7'h27}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215726.4]
  assign _T_169 = {_T_50[6:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h2,_T_50[4:0],7'h23}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215762.4]
  assign _T_200 = {_T_50[6:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h2,_T_50[4:0],7'h27}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215798.4]
  assign _T_211 = io_in[12] ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@215814.4]
  assign _T_213 = {_T_211,io_in[6:2]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215816.4]
  assign _T_219 = {_T_211,io_in[6:2],io_in[11:7],3'h0,io_in[11:7],7'h13}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215822.4]
  assign _T_228 = io_in[12] ? 10'h3ff : 10'h0; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@215836.4]
  assign _T_243 = {_T_228,io_in[8],io_in[10:9],io_in[6],io_in[7],io_in[2],io_in[11],io_in[5:3],1'h0}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215851.4]
  assign _T_306 = {_T_243[20],_T_243[10:1],_T_243[11],_T_243[19:12],5'h1,7'h6f}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215914.4]
  assign _T_321 = {_T_211,io_in[6:2],5'h0,3'h0,io_in[11:7],7'h13}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215934.4]
  assign _T_332 = |_T_213; // @[RVC.scala 91:29:freechips.rocketchip.system.DefaultRV32Config.fir@215950.4]
  assign _T_333 = _T_332 ? 7'h37 : 7'h3f; // @[RVC.scala 91:20:freechips.rocketchip.system.DefaultRV32Config.fir@215951.4]
  assign _T_336 = io_in[12] ? 15'h7fff : 15'h0; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@215954.4]
  assign _T_339 = {_T_336,io_in[6:2],12'h0}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215957.4]
  assign _T_343 = {_T_339[31:12],io_in[11:7],_T_333}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@215961.4]
  assign _T_351 = io_in[11:7] == 5'h0; // @[RVC.scala 93:14:freechips.rocketchip.system.DefaultRV32Config.fir@215974.4]
  assign _T_353 = io_in[11:7] == 5'h2; // @[RVC.scala 93:27:freechips.rocketchip.system.DefaultRV32Config.fir@215976.4]
  assign _T_354 = _T_351 | _T_353; // @[RVC.scala 93:21:freechips.rocketchip.system.DefaultRV32Config.fir@215977.4]
  assign _T_361 = _T_332 ? 7'h13 : 7'h1f; // @[RVC.scala 87:20:freechips.rocketchip.system.DefaultRV32Config.fir@215984.4]
  assign _T_364 = io_in[12] ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@215987.4]
  assign _T_379 = {_T_364,io_in[4:3],io_in[5],io_in[2],io_in[6],4'h0,io_in[11:7],3'h0,io_in[11:7],_T_361}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216002.4]
  assign _T_386_bits = _T_354 ? _T_379 : _T_343; // @[RVC.scala 93:10:freechips.rocketchip.system.DefaultRV32Config.fir@216014.4]
  assign _T_386_rd = _T_354 ? io_in[11:7] : io_in[11:7]; // @[RVC.scala 93:10:freechips.rocketchip.system.DefaultRV32Config.fir@216014.4]
  assign _T_386_rs2 = _T_354 ? _T_14 : _T_14; // @[RVC.scala 93:10:freechips.rocketchip.system.DefaultRV32Config.fir@216014.4]
  assign _T_386_rs3 = _T_354 ? io_in[31:27] : io_in[31:27]; // @[RVC.scala 93:10:freechips.rocketchip.system.DefaultRV32Config.fir@216014.4]
  assign _T_397 = {io_in[12],io_in[6:2],2'h1,io_in[9:7],3'h5,2'h1,io_in[9:7],7'h13}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216025.4]
  assign _GEN_0 = {{5'd0}, _T_397}; // @[RVC.scala 100:23:freechips.rocketchip.system.DefaultRV32Config.fir@216037.4]
  assign _T_409 = _GEN_0 | 31'h40000000; // @[RVC.scala 100:23:freechips.rocketchip.system.DefaultRV32Config.fir@216037.4]
  assign _T_422 = {_T_211,io_in[6:2],2'h1,io_in[9:7],3'h7,2'h1,io_in[9:7],7'h13}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216050.4]
  assign _T_425 = {io_in[12],io_in[6:5]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216053.4]
  assign _T_426 = _T_425 == 3'h1; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216054.4]
  assign _T_427 = _T_426 ? 3'h4 : 3'h0; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216055.4]
  assign _T_428 = _T_425 == 3'h2; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216056.4]
  assign _T_429 = _T_428 ? 3'h6 : _T_427; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216057.4]
  assign _T_430 = _T_425 == 3'h3; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216058.4]
  assign _T_431 = _T_430 ? 3'h7 : _T_429; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216059.4]
  assign _T_432 = _T_425 == 3'h4; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216060.4]
  assign _T_433 = _T_432 ? 3'h0 : _T_431; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216061.4]
  assign _T_434 = _T_425 == 3'h5; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216062.4]
  assign _T_435 = _T_434 ? 3'h0 : _T_433; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216063.4]
  assign _T_436 = _T_425 == 3'h6; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216064.4]
  assign _T_437 = _T_436 ? 3'h2 : _T_435; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216065.4]
  assign _T_438 = _T_425 == 3'h7; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216066.4]
  assign _T_439 = _T_438 ? 3'h3 : _T_437; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216067.4]
  assign _T_441 = io_in[6:5] == 2'h0; // @[RVC.scala 104:30:freechips.rocketchip.system.DefaultRV32Config.fir@216069.4]
  assign _T_442 = _T_441 ? 31'h40000000 : 31'h0; // @[RVC.scala 104:22:freechips.rocketchip.system.DefaultRV32Config.fir@216070.4]
  assign _T_444 = io_in[12] ? 7'h3b : 7'h33; // @[RVC.scala 105:22:freechips.rocketchip.system.DefaultRV32Config.fir@216072.4]
  assign _T_454 = {2'h1,io_in[4:2],2'h1,io_in[9:7],_T_439,2'h1,io_in[9:7],_T_444}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216082.4]
  assign _GEN_1 = {{6'd0}, _T_454}; // @[RVC.scala 106:43:freechips.rocketchip.system.DefaultRV32Config.fir@216083.4]
  assign _T_455 = _GEN_1 | _T_442; // @[RVC.scala 106:43:freechips.rocketchip.system.DefaultRV32Config.fir@216083.4]
  assign _T_457 = io_in[11:10] == 2'h1; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216085.4]
  assign _T_458 = _T_457 ? _T_409 : {{5'd0}, _T_397}; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216086.4]
  assign _T_459 = io_in[11:10] == 2'h2; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216087.4]
  assign _T_460 = _T_459 ? _T_422 : {{1'd0}, _T_458}; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216088.4]
  assign _T_461 = io_in[11:10] == 2'h3; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216089.4]
  assign _T_462 = _T_461 ? {{1'd0}, _T_455} : _T_460; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216090.4]
  assign _T_551 = {_T_243[20],_T_243[10:1],_T_243[11],_T_243[19:12],5'h0,7'h6f}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216184.4]
  assign _T_560 = io_in[12] ? 5'h1f : 5'h0; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultRV32Config.fir@216198.4]
  assign _T_569 = {_T_560,io_in[6:5],io_in[2],io_in[11:10],io_in[4:3],1'h0}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216207.4]
  assign _T_618 = {_T_569[12],_T_569[10:5],5'h0,2'h1,io_in[9:7],3'h0,_T_569[4:1],_T_569[11],7'h63}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216256.4]
  assign _T_685 = {_T_569[12],_T_569[10:5],5'h0,2'h1,io_in[9:7],3'h1,_T_569[4:1],_T_569[11],7'h63}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216328.4]
  assign _T_691 = |io_in[11:7]; // @[RVC.scala 114:27:freechips.rocketchip.system.DefaultRV32Config.fir@216339.4]
  assign _T_692 = _T_691 ? 7'h3 : 7'h1f; // @[RVC.scala 114:23:freechips.rocketchip.system.DefaultRV32Config.fir@216340.4]
  assign _T_701 = {io_in[12],io_in[6:2],io_in[11:7],3'h1,io_in[11:7],7'h13}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216349.4]
  assign _T_717 = {io_in[4:2],io_in[12],io_in[6:5],3'h0,5'h2,3'h3,io_in[11:7],7'h7}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216370.4]
  assign _T_732 = {io_in[3:2],io_in[12],io_in[6:4],2'h0,5'h2,3'h2,io_in[11:7],_T_692}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216390.4]
  assign _T_747 = {io_in[3:2],io_in[12],io_in[6:4],2'h0,5'h2,3'h2,io_in[11:7],7'h7}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216410.4]
  assign _T_757 = {io_in[6:2],5'h0,3'h0,io_in[11:7],7'h33}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216425.4]
  assign _T_768 = {io_in[6:2],io_in[11:7],3'h0,io_in[11:7],7'h33}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216441.4]
  assign _T_779 = {io_in[6:2],io_in[11:7],3'h0,12'h67}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216457.4]
  assign _T_781 = {_T_779[24:7],7'h1f}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216459.4]
  assign _T_784 = _T_691 ? _T_779 : _T_781; // @[RVC.scala 135:33:freechips.rocketchip.system.DefaultRV32Config.fir@216462.4]
  assign _T_790 = |io_in[6:2]; // @[RVC.scala 136:27:freechips.rocketchip.system.DefaultRV32Config.fir@216473.4]
  assign _T_761_bits = {{7'd0}, _T_757}; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@216429.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@216430.4]
  assign _T_788_bits = {{7'd0}, _T_784}; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@216466.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@216467.4]
  assign _T_791_bits = _T_790 ? _T_761_bits : _T_788_bits; // @[RVC.scala 136:22:freechips.rocketchip.system.DefaultRV32Config.fir@216474.4]
  assign _T_791_rd = _T_790 ? io_in[11:7] : 5'h0; // @[RVC.scala 136:22:freechips.rocketchip.system.DefaultRV32Config.fir@216474.4]
  assign _T_791_rs1 = _T_790 ? 5'h0 : io_in[11:7]; // @[RVC.scala 136:22:freechips.rocketchip.system.DefaultRV32Config.fir@216474.4]
  assign _T_791_rs2 = _T_790 ? io_in[6:2] : io_in[6:2]; // @[RVC.scala 136:22:freechips.rocketchip.system.DefaultRV32Config.fir@216474.4]
  assign _T_791_rs3 = _T_790 ? io_in[31:27] : io_in[31:27]; // @[RVC.scala 136:22:freechips.rocketchip.system.DefaultRV32Config.fir@216474.4]
  assign _T_797 = {io_in[6:2],io_in[11:7],3'h0,12'he7}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216480.4]
  assign _T_799 = {_T_779[24:7],7'h73}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216482.4]
  assign _T_800 = _T_799 | 25'h100000; // @[RVC.scala 138:46:freechips.rocketchip.system.DefaultRV32Config.fir@216483.4]
  assign _T_803 = _T_691 ? _T_797 : _T_800; // @[RVC.scala 139:33:freechips.rocketchip.system.DefaultRV32Config.fir@216486.4]
  assign _T_773_bits = {{7'd0}, _T_768}; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@216446.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@216447.4]
  assign _T_807_bits = {{7'd0}, _T_803}; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@216490.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@216491.4]
  assign _T_810_bits = _T_790 ? _T_773_bits : _T_807_bits; // @[RVC.scala 140:25:freechips.rocketchip.system.DefaultRV32Config.fir@216498.4]
  assign _T_810_rd = _T_790 ? io_in[11:7] : 5'h1; // @[RVC.scala 140:25:freechips.rocketchip.system.DefaultRV32Config.fir@216498.4]
  assign _T_810_rs1 = _T_790 ? io_in[11:7] : io_in[11:7]; // @[RVC.scala 140:25:freechips.rocketchip.system.DefaultRV32Config.fir@216498.4]
  assign _T_812_bits = io_in[12] ? _T_810_bits : _T_791_bits; // @[RVC.scala 141:10:freechips.rocketchip.system.DefaultRV32Config.fir@216500.4]
  assign _T_812_rd = io_in[12] ? _T_810_rd : _T_791_rd; // @[RVC.scala 141:10:freechips.rocketchip.system.DefaultRV32Config.fir@216500.4]
  assign _T_812_rs1 = io_in[12] ? _T_810_rs1 : _T_791_rs1; // @[RVC.scala 141:10:freechips.rocketchip.system.DefaultRV32Config.fir@216500.4]
  assign _T_812_rs2 = io_in[12] ? _T_791_rs2 : _T_791_rs2; // @[RVC.scala 141:10:freechips.rocketchip.system.DefaultRV32Config.fir@216500.4]
  assign _T_812_rs3 = io_in[12] ? _T_791_rs3 : _T_791_rs3; // @[RVC.scala 141:10:freechips.rocketchip.system.DefaultRV32Config.fir@216500.4]
  assign _T_816 = {io_in[9:7],io_in[12:10],3'h0}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216504.4]
  assign _T_828 = {_T_816[8:5],io_in[6:2],5'h2,3'h3,_T_816[4:0],7'h27}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216516.4]
  assign _T_836 = {io_in[8:7],io_in[12:9],2'h0}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216529.4]
  assign _T_848 = {_T_836[7:5],io_in[6:2],5'h2,3'h2,_T_836[4:0],7'h23}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216541.4]
  assign _T_868 = {_T_836[7:5],io_in[6:2],5'h2,3'h2,_T_836[4:0],7'h27}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216566.4]
  assign _T_915 = {io_in[1:0],io_in[15:13]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@216658.4]
  assign _T_916 = _T_915 == 5'h1; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216659.4]
  assign _T_44_bits = {{4'd0}, _T_36}; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@215612.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@215613.4]
  assign _T_24_bits = {{2'd0}, _T_18}; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@215587.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@215588.4]
  assign _T_917_bits = _T_916 ? _T_44_bits : _T_24_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216660.4]
  assign _T_917_rd = _T_916 ? _T_14 : _T_14; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216660.4]
  assign _T_917_rs1 = _T_916 ? _T_30 : 5'h2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216660.4]
  assign _T_917_rs3 = _T_916 ? io_in[31:27] : io_in[31:27]; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216660.4]
  assign _T_918 = _T_915 == 5'h2; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216661.4]
  assign _T_66_bits = {{5'd0}, _T_58}; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@215639.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@215640.4]
  assign _T_919_bits = _T_918 ? _T_66_bits : _T_917_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216662.4]
  assign _T_919_rd = _T_918 ? _T_14 : _T_917_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216662.4]
  assign _T_919_rs1 = _T_918 ? _T_30 : _T_917_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216662.4]
  assign _T_919_rs3 = _T_918 ? io_in[31:27] : _T_917_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216662.4]
  assign _T_920 = _T_915 == 5'h3; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216663.4]
  assign _T_88_bits = {{5'd0}, _T_80}; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@215666.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@215667.4]
  assign _T_921_bits = _T_920 ? _T_88_bits : _T_919_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216664.4]
  assign _T_921_rd = _T_920 ? _T_14 : _T_919_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216664.4]
  assign _T_921_rs1 = _T_920 ? _T_30 : _T_919_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216664.4]
  assign _T_921_rs3 = _T_920 ? io_in[31:27] : _T_919_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216664.4]
  assign _T_922 = _T_915 == 5'h4; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216665.4]
  assign _T_119_bits = {{5'd0}, _T_111}; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@215702.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@215703.4]
  assign _T_923_bits = _T_922 ? _T_119_bits : _T_921_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216666.4]
  assign _T_923_rd = _T_922 ? _T_14 : _T_921_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216666.4]
  assign _T_923_rs1 = _T_922 ? _T_30 : _T_921_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216666.4]
  assign _T_923_rs3 = _T_922 ? io_in[31:27] : _T_921_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216666.4]
  assign _T_924 = _T_915 == 5'h5; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216667.4]
  assign _T_146_bits = {{4'd0}, _T_138}; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@215734.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@215735.4]
  assign _T_925_bits = _T_924 ? _T_146_bits : _T_923_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216668.4]
  assign _T_925_rd = _T_924 ? _T_14 : _T_923_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216668.4]
  assign _T_925_rs1 = _T_924 ? _T_30 : _T_923_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216668.4]
  assign _T_925_rs3 = _T_924 ? io_in[31:27] : _T_923_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216668.4]
  assign _T_926 = _T_915 == 5'h6; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216669.4]
  assign _T_177_bits = {{5'd0}, _T_169}; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@215770.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@215771.4]
  assign _T_927_bits = _T_926 ? _T_177_bits : _T_925_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216670.4]
  assign _T_927_rd = _T_926 ? _T_14 : _T_925_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216670.4]
  assign _T_927_rs1 = _T_926 ? _T_30 : _T_925_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216670.4]
  assign _T_927_rs3 = _T_926 ? io_in[31:27] : _T_925_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216670.4]
  assign _T_928 = _T_915 == 5'h7; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216671.4]
  assign _T_208_bits = {{5'd0}, _T_200}; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@215806.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@215807.4]
  assign _T_929_bits = _T_928 ? _T_208_bits : _T_927_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216672.4]
  assign _T_929_rd = _T_928 ? _T_14 : _T_927_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216672.4]
  assign _T_929_rs1 = _T_928 ? _T_30 : _T_927_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216672.4]
  assign _T_929_rs3 = _T_928 ? io_in[31:27] : _T_927_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216672.4]
  assign _T_930 = _T_915 == 5'h8; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216673.4]
  assign _T_931_bits = _T_930 ? _T_219 : _T_929_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216674.4]
  assign _T_931_rd = _T_930 ? io_in[11:7] : _T_929_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216674.4]
  assign _T_931_rs1 = _T_930 ? io_in[11:7] : _T_929_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216674.4]
  assign _T_931_rs2 = _T_930 ? _T_14 : _T_929_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216674.4]
  assign _T_931_rs3 = _T_930 ? io_in[31:27] : _T_929_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216674.4]
  assign _T_932 = _T_915 == 5'h9; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216675.4]
  assign _T_933_bits = _T_932 ? _T_306 : _T_931_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216676.4]
  assign _T_933_rd = _T_932 ? 5'h1 : _T_931_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216676.4]
  assign _T_933_rs1 = _T_932 ? io_in[11:7] : _T_931_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216676.4]
  assign _T_933_rs2 = _T_932 ? _T_14 : _T_931_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216676.4]
  assign _T_933_rs3 = _T_932 ? io_in[31:27] : _T_931_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216676.4]
  assign _T_934 = _T_915 == 5'ha; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216677.4]
  assign _T_935_bits = _T_934 ? _T_321 : _T_933_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216678.4]
  assign _T_935_rd = _T_934 ? io_in[11:7] : _T_933_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216678.4]
  assign _T_935_rs1 = _T_934 ? 5'h0 : _T_933_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216678.4]
  assign _T_935_rs2 = _T_934 ? _T_14 : _T_933_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216678.4]
  assign _T_935_rs3 = _T_934 ? io_in[31:27] : _T_933_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216678.4]
  assign _T_936 = _T_915 == 5'hb; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216679.4]
  assign _T_937_bits = _T_936 ? _T_386_bits : _T_935_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216680.4]
  assign _T_937_rd = _T_936 ? _T_386_rd : _T_935_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216680.4]
  assign _T_937_rs1 = _T_936 ? _T_386_rd : _T_935_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216680.4]
  assign _T_937_rs2 = _T_936 ? _T_386_rs2 : _T_935_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216680.4]
  assign _T_937_rs3 = _T_936 ? _T_386_rs3 : _T_935_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216680.4]
  assign _T_938 = _T_915 == 5'hc; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216681.4]
  assign _T_939_bits = _T_938 ? _T_462 : _T_937_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216682.4]
  assign _T_939_rd = _T_938 ? _T_30 : _T_937_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216682.4]
  assign _T_939_rs1 = _T_938 ? _T_30 : _T_937_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216682.4]
  assign _T_939_rs2 = _T_938 ? _T_14 : _T_937_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216682.4]
  assign _T_939_rs3 = _T_938 ? io_in[31:27] : _T_937_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216682.4]
  assign _T_940 = _T_915 == 5'hd; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216683.4]
  assign _T_941_bits = _T_940 ? _T_551 : _T_939_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216684.4]
  assign _T_941_rd = _T_940 ? 5'h0 : _T_939_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216684.4]
  assign _T_941_rs1 = _T_940 ? _T_30 : _T_939_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216684.4]
  assign _T_941_rs2 = _T_940 ? _T_14 : _T_939_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216684.4]
  assign _T_941_rs3 = _T_940 ? io_in[31:27] : _T_939_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216684.4]
  assign _T_942 = _T_915 == 5'he; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216685.4]
  assign _T_943_bits = _T_942 ? _T_618 : _T_941_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216686.4]
  assign _T_943_rd = _T_942 ? _T_30 : _T_941_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216686.4]
  assign _T_943_rs1 = _T_942 ? _T_30 : _T_941_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216686.4]
  assign _T_943_rs2 = _T_942 ? 5'h0 : _T_941_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216686.4]
  assign _T_943_rs3 = _T_942 ? io_in[31:27] : _T_941_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216686.4]
  assign _T_944 = _T_915 == 5'hf; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216687.4]
  assign _T_945_bits = _T_944 ? _T_685 : _T_943_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216688.4]
  assign _T_945_rd = _T_944 ? 5'h0 : _T_943_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216688.4]
  assign _T_945_rs1 = _T_944 ? _T_30 : _T_943_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216688.4]
  assign _T_945_rs2 = _T_944 ? 5'h0 : _T_943_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216688.4]
  assign _T_945_rs3 = _T_944 ? io_in[31:27] : _T_943_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216688.4]
  assign _T_946 = _T_915 == 5'h10; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216689.4]
  assign _T_706_bits = {{6'd0}, _T_701}; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@216354.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@216355.4]
  assign _T_947_bits = _T_946 ? _T_706_bits : _T_945_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216690.4]
  assign _T_947_rd = _T_946 ? io_in[11:7] : _T_945_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216690.4]
  assign _T_947_rs1 = _T_946 ? io_in[11:7] : _T_945_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216690.4]
  assign _T_947_rs2 = _T_946 ? io_in[6:2] : _T_945_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216690.4]
  assign _T_947_rs3 = _T_946 ? io_in[31:27] : _T_945_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216690.4]
  assign _T_948 = _T_915 == 5'h11; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216691.4]
  assign _T_721_bits = {{3'd0}, _T_717}; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@216374.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@216375.4]
  assign _T_949_bits = _T_948 ? _T_721_bits : _T_947_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216692.4]
  assign _T_949_rd = _T_948 ? io_in[11:7] : _T_947_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216692.4]
  assign _T_949_rs1 = _T_948 ? 5'h2 : _T_947_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216692.4]
  assign _T_949_rs2 = _T_948 ? io_in[6:2] : _T_947_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216692.4]
  assign _T_949_rs3 = _T_948 ? io_in[31:27] : _T_947_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216692.4]
  assign _T_950 = _T_915 == 5'h12; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216693.4]
  assign _T_736_bits = {{4'd0}, _T_732}; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@216394.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@216395.4]
  assign _T_951_bits = _T_950 ? _T_736_bits : _T_949_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216694.4]
  assign _T_951_rd = _T_950 ? io_in[11:7] : _T_949_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216694.4]
  assign _T_951_rs1 = _T_950 ? 5'h2 : _T_949_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216694.4]
  assign _T_951_rs2 = _T_950 ? io_in[6:2] : _T_949_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216694.4]
  assign _T_951_rs3 = _T_950 ? io_in[31:27] : _T_949_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216694.4]
  assign _T_952 = _T_915 == 5'h13; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216695.4]
  assign _T_751_bits = {{4'd0}, _T_747}; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@216414.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@216415.4]
  assign _T_953_bits = _T_952 ? _T_751_bits : _T_951_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216696.4]
  assign _T_953_rd = _T_952 ? io_in[11:7] : _T_951_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216696.4]
  assign _T_953_rs1 = _T_952 ? 5'h2 : _T_951_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216696.4]
  assign _T_953_rs2 = _T_952 ? io_in[6:2] : _T_951_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216696.4]
  assign _T_953_rs3 = _T_952 ? io_in[31:27] : _T_951_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216696.4]
  assign _T_954 = _T_915 == 5'h14; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216697.4]
  assign _T_955_bits = _T_954 ? _T_812_bits : _T_953_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216698.4]
  assign _T_955_rd = _T_954 ? _T_812_rd : _T_953_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216698.4]
  assign _T_955_rs1 = _T_954 ? _T_812_rs1 : _T_953_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216698.4]
  assign _T_955_rs2 = _T_954 ? _T_812_rs2 : _T_953_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216698.4]
  assign _T_955_rs3 = _T_954 ? _T_812_rs3 : _T_953_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216698.4]
  assign _T_956 = _T_915 == 5'h15; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216699.4]
  assign _T_832_bits = {{3'd0}, _T_828}; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@216520.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@216521.4]
  assign _T_957_bits = _T_956 ? _T_832_bits : _T_955_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216700.4]
  assign _T_957_rd = _T_956 ? io_in[11:7] : _T_955_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216700.4]
  assign _T_957_rs1 = _T_956 ? 5'h2 : _T_955_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216700.4]
  assign _T_957_rs2 = _T_956 ? io_in[6:2] : _T_955_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216700.4]
  assign _T_957_rs3 = _T_956 ? io_in[31:27] : _T_955_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216700.4]
  assign _T_958 = _T_915 == 5'h16; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216701.4]
  assign _T_852_bits = {{4'd0}, _T_848}; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@216545.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@216546.4]
  assign _T_959_bits = _T_958 ? _T_852_bits : _T_957_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216702.4]
  assign _T_959_rd = _T_958 ? io_in[11:7] : _T_957_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216702.4]
  assign _T_959_rs1 = _T_958 ? 5'h2 : _T_957_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216702.4]
  assign _T_959_rs2 = _T_958 ? io_in[6:2] : _T_957_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216702.4]
  assign _T_959_rs3 = _T_958 ? io_in[31:27] : _T_957_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216702.4]
  assign _T_960 = _T_915 == 5'h17; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216703.4]
  assign _T_872_bits = {{4'd0}, _T_868}; // @[RVC.scala 22:19:freechips.rocketchip.system.DefaultRV32Config.fir@216570.4 RVC.scala 23:14:freechips.rocketchip.system.DefaultRV32Config.fir@216571.4]
  assign _T_961_bits = _T_960 ? _T_872_bits : _T_959_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216704.4]
  assign _T_961_rd = _T_960 ? io_in[11:7] : _T_959_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216704.4]
  assign _T_961_rs1 = _T_960 ? 5'h2 : _T_959_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216704.4]
  assign _T_961_rs2 = _T_960 ? io_in[6:2] : _T_959_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216704.4]
  assign _T_961_rs3 = _T_960 ? io_in[31:27] : _T_959_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216704.4]
  assign _T_962 = _T_915 == 5'h18; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216705.4]
  assign _T_963_bits = _T_962 ? io_in : _T_961_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216706.4]
  assign _T_963_rd = _T_962 ? io_in[11:7] : _T_961_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216706.4]
  assign _T_963_rs1 = _T_962 ? io_in[19:15] : _T_961_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216706.4]
  assign _T_963_rs2 = _T_962 ? io_in[24:20] : _T_961_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216706.4]
  assign _T_963_rs3 = _T_962 ? io_in[31:27] : _T_961_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216706.4]
  assign _T_964 = _T_915 == 5'h19; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216707.4]
  assign _T_965_bits = _T_964 ? io_in : _T_963_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216708.4]
  assign _T_965_rd = _T_964 ? io_in[11:7] : _T_963_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216708.4]
  assign _T_965_rs1 = _T_964 ? io_in[19:15] : _T_963_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216708.4]
  assign _T_965_rs2 = _T_964 ? io_in[24:20] : _T_963_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216708.4]
  assign _T_965_rs3 = _T_964 ? io_in[31:27] : _T_963_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216708.4]
  assign _T_966 = _T_915 == 5'h1a; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216709.4]
  assign _T_967_bits = _T_966 ? io_in : _T_965_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216710.4]
  assign _T_967_rd = _T_966 ? io_in[11:7] : _T_965_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216710.4]
  assign _T_967_rs1 = _T_966 ? io_in[19:15] : _T_965_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216710.4]
  assign _T_967_rs2 = _T_966 ? io_in[24:20] : _T_965_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216710.4]
  assign _T_967_rs3 = _T_966 ? io_in[31:27] : _T_965_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216710.4]
  assign _T_968 = _T_915 == 5'h1b; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216711.4]
  assign _T_969_bits = _T_968 ? io_in : _T_967_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216712.4]
  assign _T_969_rd = _T_968 ? io_in[11:7] : _T_967_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216712.4]
  assign _T_969_rs1 = _T_968 ? io_in[19:15] : _T_967_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216712.4]
  assign _T_969_rs2 = _T_968 ? io_in[24:20] : _T_967_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216712.4]
  assign _T_969_rs3 = _T_968 ? io_in[31:27] : _T_967_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216712.4]
  assign _T_970 = _T_915 == 5'h1c; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216713.4]
  assign _T_971_bits = _T_970 ? io_in : _T_969_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216714.4]
  assign _T_971_rd = _T_970 ? io_in[11:7] : _T_969_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216714.4]
  assign _T_971_rs1 = _T_970 ? io_in[19:15] : _T_969_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216714.4]
  assign _T_971_rs2 = _T_970 ? io_in[24:20] : _T_969_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216714.4]
  assign _T_971_rs3 = _T_970 ? io_in[31:27] : _T_969_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216714.4]
  assign _T_972 = _T_915 == 5'h1d; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216715.4]
  assign _T_973_bits = _T_972 ? io_in : _T_971_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216716.4]
  assign _T_973_rd = _T_972 ? io_in[11:7] : _T_971_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216716.4]
  assign _T_973_rs1 = _T_972 ? io_in[19:15] : _T_971_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216716.4]
  assign _T_973_rs2 = _T_972 ? io_in[24:20] : _T_971_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216716.4]
  assign _T_973_rs3 = _T_972 ? io_in[31:27] : _T_971_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216716.4]
  assign _T_974 = _T_915 == 5'h1e; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216717.4]
  assign _T_975_bits = _T_974 ? io_in : _T_973_bits; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216718.4]
  assign _T_975_rd = _T_974 ? io_in[11:7] : _T_973_rd; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216718.4]
  assign _T_975_rs1 = _T_974 ? io_in[19:15] : _T_973_rs1; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216718.4]
  assign _T_975_rs2 = _T_974 ? io_in[24:20] : _T_973_rs2; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216718.4]
  assign _T_975_rs3 = _T_974 ? io_in[31:27] : _T_973_rs3; // @[package.scala 32:76:freechips.rocketchip.system.DefaultRV32Config.fir@216718.4]
  assign _T_976 = _T_915 == 5'h1f; // @[package.scala 32:86:freechips.rocketchip.system.DefaultRV32Config.fir@216719.4]
  assign io_out_bits = _T_976 ? io_in : _T_975_bits; // @[RVC.scala 165:12:freechips.rocketchip.system.DefaultRV32Config.fir@216725.4]
  assign io_out_rd = _T_976 ? io_in[11:7] : _T_975_rd; // @[RVC.scala 165:12:freechips.rocketchip.system.DefaultRV32Config.fir@216724.4]
  assign io_out_rs1 = _T_976 ? io_in[19:15] : _T_975_rs1; // @[RVC.scala 165:12:freechips.rocketchip.system.DefaultRV32Config.fir@216723.4]
  assign io_out_rs2 = _T_976 ? io_in[24:20] : _T_975_rs2; // @[RVC.scala 165:12:freechips.rocketchip.system.DefaultRV32Config.fir@216722.4]
  assign io_out_rs3 = _T_976 ? io_in[31:27] : _T_975_rs3; // @[RVC.scala 165:12:freechips.rocketchip.system.DefaultRV32Config.fir@216721.4]
  assign io_rvc = io_in[1:0] != 2'h3; // @[RVC.scala 164:12:freechips.rocketchip.system.DefaultRV32Config.fir@215564.4]
endmodule
