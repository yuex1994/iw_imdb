module IntSyncSyncCrossingSink_1( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@210973.2]
  input   auto_in_sync_0, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@210976.4]
  output  auto_out_0 // @[:freechips.rocketchip.system.DefaultRV32Config.fir@210976.4]
);
  assign auto_out_0 = auto_in_sync_0; // @[LazyModule.scala 305:12:freechips.rocketchip.system.DefaultRV32Config.fir@210985.4]
endmodule
