module BreakpointUnit( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@224124.2]
  input         io_status_debug, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@224127.4]
  input  [1:0]  io_status_prv, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@224127.4]
  input         io_bp_0_control_action, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@224127.4]
  input  [1:0]  io_bp_0_control_tmatch, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@224127.4]
  input         io_bp_0_control_m, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@224127.4]
  input         io_bp_0_control_s, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@224127.4]
  input         io_bp_0_control_u, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@224127.4]
  input         io_bp_0_control_x, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@224127.4]
  input         io_bp_0_control_w, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@224127.4]
  input         io_bp_0_control_r, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@224127.4]
  input  [31:0] io_bp_0_address, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@224127.4]
  input  [31:0] io_pc, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@224127.4]
  input  [31:0] io_ea, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@224127.4]
  output        io_xcpt_if, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@224127.4]
  output        io_xcpt_ld, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@224127.4]
  output        io_xcpt_st, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@224127.4]
  output        io_debug_if, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@224127.4]
  output        io_debug_ld, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@224127.4]
  output        io_debug_st // @[:freechips.rocketchip.system.DefaultRV32Config.fir@224127.4]
);
  wire  _T; // @[Breakpoint.scala 31:35:freechips.rocketchip.system.DefaultRV32Config.fir@224135.4]
  wire [3:0] _T_3; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@224138.4]
  wire [3:0] _T_4; // @[Breakpoint.scala 31:68:freechips.rocketchip.system.DefaultRV32Config.fir@224139.4]
  wire  _T_6; // @[Breakpoint.scala 31:50:freechips.rocketchip.system.DefaultRV32Config.fir@224141.4]
  wire  _T_7; // @[Breakpoint.scala 83:16:freechips.rocketchip.system.DefaultRV32Config.fir@224142.4]
  wire  _T_9; // @[Breakpoint.scala 45:8:freechips.rocketchip.system.DefaultRV32Config.fir@224144.4]
  wire  _T_11; // @[Breakpoint.scala 45:20:freechips.rocketchip.system.DefaultRV32Config.fir@224146.4]
  wire [31:0] _T_12; // @[Breakpoint.scala 42:6:freechips.rocketchip.system.DefaultRV32Config.fir@224147.4]
  wire  _T_15; // @[Breakpoint.scala 39:73:freechips.rocketchip.system.DefaultRV32Config.fir@224150.4]
  wire  _T_17; // @[Breakpoint.scala 39:73:freechips.rocketchip.system.DefaultRV32Config.fir@224152.4]
  wire  _T_19; // @[Breakpoint.scala 39:73:freechips.rocketchip.system.DefaultRV32Config.fir@224154.4]
  wire [3:0] _T_22; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@224157.4]
  wire [31:0] _GEN_11; // @[Breakpoint.scala 42:9:freechips.rocketchip.system.DefaultRV32Config.fir@224158.4]
  wire [31:0] _T_23; // @[Breakpoint.scala 42:9:freechips.rocketchip.system.DefaultRV32Config.fir@224158.4]
  wire [31:0] _T_24; // @[Breakpoint.scala 42:24:freechips.rocketchip.system.DefaultRV32Config.fir@224159.4]
  wire [31:0] _T_35; // @[Breakpoint.scala 42:33:freechips.rocketchip.system.DefaultRV32Config.fir@224170.4]
  wire  _T_36; // @[Breakpoint.scala 42:19:freechips.rocketchip.system.DefaultRV32Config.fir@224171.4]
  wire  _T_37; // @[Breakpoint.scala 48:8:freechips.rocketchip.system.DefaultRV32Config.fir@224172.4]
  wire  _T_38; // @[Breakpoint.scala 83:32:freechips.rocketchip.system.DefaultRV32Config.fir@224173.4]
  wire  _T_39; // @[Breakpoint.scala 84:16:freechips.rocketchip.system.DefaultRV32Config.fir@224174.4]
  wire  _T_70; // @[Breakpoint.scala 84:32:freechips.rocketchip.system.DefaultRV32Config.fir@224205.4]
  wire  _T_71; // @[Breakpoint.scala 85:16:freechips.rocketchip.system.DefaultRV32Config.fir@224206.4]
  wire  _T_73; // @[Breakpoint.scala 45:8:freechips.rocketchip.system.DefaultRV32Config.fir@224208.4]
  wire  _T_75; // @[Breakpoint.scala 45:20:freechips.rocketchip.system.DefaultRV32Config.fir@224210.4]
  wire [31:0] _T_76; // @[Breakpoint.scala 42:6:freechips.rocketchip.system.DefaultRV32Config.fir@224211.4]
  wire [31:0] _T_87; // @[Breakpoint.scala 42:9:freechips.rocketchip.system.DefaultRV32Config.fir@224222.4]
  wire  _T_100; // @[Breakpoint.scala 42:19:freechips.rocketchip.system.DefaultRV32Config.fir@224235.4]
  wire  _T_101; // @[Breakpoint.scala 48:8:freechips.rocketchip.system.DefaultRV32Config.fir@224236.4]
  wire  _T_102; // @[Breakpoint.scala 85:32:freechips.rocketchip.system.DefaultRV32Config.fir@224237.4]
  wire  _T_106; // @[Breakpoint.scala 95:51:freechips.rocketchip.system.DefaultRV32Config.fir@224247.6]
  assign _T = ~io_status_debug; // @[Breakpoint.scala 31:35:freechips.rocketchip.system.DefaultRV32Config.fir@224135.4]
  assign _T_3 = {io_bp_0_control_m,1'h0,io_bp_0_control_s,io_bp_0_control_u}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@224138.4]
  assign _T_4 = _T_3 >> io_status_prv; // @[Breakpoint.scala 31:68:freechips.rocketchip.system.DefaultRV32Config.fir@224139.4]
  assign _T_6 = _T & _T_4[0]; // @[Breakpoint.scala 31:50:freechips.rocketchip.system.DefaultRV32Config.fir@224141.4]
  assign _T_7 = _T_6 & io_bp_0_control_r; // @[Breakpoint.scala 83:16:freechips.rocketchip.system.DefaultRV32Config.fir@224142.4]
  assign _T_9 = io_ea >= io_bp_0_address; // @[Breakpoint.scala 45:8:freechips.rocketchip.system.DefaultRV32Config.fir@224144.4]
  assign _T_11 = _T_9 ^ io_bp_0_control_tmatch[0]; // @[Breakpoint.scala 45:20:freechips.rocketchip.system.DefaultRV32Config.fir@224146.4]
  assign _T_12 = ~io_ea; // @[Breakpoint.scala 42:6:freechips.rocketchip.system.DefaultRV32Config.fir@224147.4]
  assign _T_15 = io_bp_0_control_tmatch[0] & io_bp_0_address[0]; // @[Breakpoint.scala 39:73:freechips.rocketchip.system.DefaultRV32Config.fir@224150.4]
  assign _T_17 = _T_15 & io_bp_0_address[1]; // @[Breakpoint.scala 39:73:freechips.rocketchip.system.DefaultRV32Config.fir@224152.4]
  assign _T_19 = _T_17 & io_bp_0_address[2]; // @[Breakpoint.scala 39:73:freechips.rocketchip.system.DefaultRV32Config.fir@224154.4]
  assign _T_22 = {_T_19,_T_17,_T_15,io_bp_0_control_tmatch[0]}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@224157.4]
  assign _GEN_11 = {{28'd0}, _T_22}; // @[Breakpoint.scala 42:9:freechips.rocketchip.system.DefaultRV32Config.fir@224158.4]
  assign _T_23 = _T_12 | _GEN_11; // @[Breakpoint.scala 42:9:freechips.rocketchip.system.DefaultRV32Config.fir@224158.4]
  assign _T_24 = ~io_bp_0_address; // @[Breakpoint.scala 42:24:freechips.rocketchip.system.DefaultRV32Config.fir@224159.4]
  assign _T_35 = _T_24 | _GEN_11; // @[Breakpoint.scala 42:33:freechips.rocketchip.system.DefaultRV32Config.fir@224170.4]
  assign _T_36 = _T_23 == _T_35; // @[Breakpoint.scala 42:19:freechips.rocketchip.system.DefaultRV32Config.fir@224171.4]
  assign _T_37 = io_bp_0_control_tmatch[1] ? _T_11 : _T_36; // @[Breakpoint.scala 48:8:freechips.rocketchip.system.DefaultRV32Config.fir@224172.4]
  assign _T_38 = _T_7 & _T_37; // @[Breakpoint.scala 83:32:freechips.rocketchip.system.DefaultRV32Config.fir@224173.4]
  assign _T_39 = _T_6 & io_bp_0_control_w; // @[Breakpoint.scala 84:16:freechips.rocketchip.system.DefaultRV32Config.fir@224174.4]
  assign _T_70 = _T_39 & _T_37; // @[Breakpoint.scala 84:32:freechips.rocketchip.system.DefaultRV32Config.fir@224205.4]
  assign _T_71 = _T_6 & io_bp_0_control_x; // @[Breakpoint.scala 85:16:freechips.rocketchip.system.DefaultRV32Config.fir@224206.4]
  assign _T_73 = io_pc >= io_bp_0_address; // @[Breakpoint.scala 45:8:freechips.rocketchip.system.DefaultRV32Config.fir@224208.4]
  assign _T_75 = _T_73 ^ io_bp_0_control_tmatch[0]; // @[Breakpoint.scala 45:20:freechips.rocketchip.system.DefaultRV32Config.fir@224210.4]
  assign _T_76 = ~io_pc; // @[Breakpoint.scala 42:6:freechips.rocketchip.system.DefaultRV32Config.fir@224211.4]
  assign _T_87 = _T_76 | _GEN_11; // @[Breakpoint.scala 42:9:freechips.rocketchip.system.DefaultRV32Config.fir@224222.4]
  assign _T_100 = _T_87 == _T_35; // @[Breakpoint.scala 42:19:freechips.rocketchip.system.DefaultRV32Config.fir@224235.4]
  assign _T_101 = io_bp_0_control_tmatch[1] ? _T_75 : _T_100; // @[Breakpoint.scala 48:8:freechips.rocketchip.system.DefaultRV32Config.fir@224236.4]
  assign _T_102 = _T_71 & _T_101; // @[Breakpoint.scala 85:32:freechips.rocketchip.system.DefaultRV32Config.fir@224237.4]
  assign _T_106 = ~io_bp_0_control_action; // @[Breakpoint.scala 95:51:freechips.rocketchip.system.DefaultRV32Config.fir@224247.6]
  assign io_xcpt_if = _T_102 & _T_106; // @[Breakpoint.scala 74:14:freechips.rocketchip.system.DefaultRV32Config.fir@224129.4 Breakpoint.scala 97:40:freechips.rocketchip.system.DefaultRV32Config.fir@224268.6]
  assign io_xcpt_ld = _T_38 & _T_106; // @[Breakpoint.scala 75:14:freechips.rocketchip.system.DefaultRV32Config.fir@224130.4 Breakpoint.scala 95:40:freechips.rocketchip.system.DefaultRV32Config.fir@224248.6]
  assign io_xcpt_st = _T_70 & _T_106; // @[Breakpoint.scala 76:14:freechips.rocketchip.system.DefaultRV32Config.fir@224131.4 Breakpoint.scala 96:40:freechips.rocketchip.system.DefaultRV32Config.fir@224258.6]
  assign io_debug_if = _T_102 & io_bp_0_control_action; // @[Breakpoint.scala 77:15:freechips.rocketchip.system.DefaultRV32Config.fir@224132.4 Breakpoint.scala 97:73:freechips.rocketchip.system.DefaultRV32Config.fir@224270.6]
  assign io_debug_ld = _T_38 & io_bp_0_control_action; // @[Breakpoint.scala 78:15:freechips.rocketchip.system.DefaultRV32Config.fir@224133.4 Breakpoint.scala 95:73:freechips.rocketchip.system.DefaultRV32Config.fir@224250.6]
  assign io_debug_st = _T_70 & io_bp_0_control_action; // @[Breakpoint.scala 79:15:freechips.rocketchip.system.DefaultRV32Config.fir@224134.4 Breakpoint.scala 96:73:freechips.rocketchip.system.DefaultRV32Config.fir@224260.6]
endmodule
