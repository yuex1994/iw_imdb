module ALU( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@223130.2]
  input  [3:0]  io_fn, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@223133.4]
  input  [31:0] io_in2, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@223133.4]
  input  [31:0] io_in1, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@223133.4]
  output [31:0] io_out, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@223133.4]
  output [31:0] io_adder_out, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@223133.4]
  output        io_cmp_out // @[:freechips.rocketchip.system.DefaultRV32Config.fir@223133.4]
);
  wire [31:0] _T_1; // @[ALU.scala 62:35:freechips.rocketchip.system.DefaultRV32Config.fir@223139.4]
  wire [31:0] in2_inv; // @[ALU.scala 62:20:freechips.rocketchip.system.DefaultRV32Config.fir@223140.4]
  wire [31:0] in1_xor_in2; // @[ALU.scala 63:28:freechips.rocketchip.system.DefaultRV32Config.fir@223141.4]
  wire [31:0] _T_3; // @[ALU.scala 64:26:freechips.rocketchip.system.DefaultRV32Config.fir@223143.4]
  wire [31:0] _GEN_0; // @[ALU.scala 64:36:freechips.rocketchip.system.DefaultRV32Config.fir@223145.4]
  wire  _T_9; // @[ALU.scala 68:24:freechips.rocketchip.system.DefaultRV32Config.fir@223150.4]
  wire  _T_14; // @[ALU.scala 69:8:freechips.rocketchip.system.DefaultRV32Config.fir@223155.4]
  wire  slt; // @[ALU.scala 68:8:freechips.rocketchip.system.DefaultRV32Config.fir@223156.4]
  wire  _T_17; // @[ALU.scala 44:26:freechips.rocketchip.system.DefaultRV32Config.fir@223159.4]
  wire  _T_18; // @[ALU.scala 70:68:freechips.rocketchip.system.DefaultRV32Config.fir@223160.4]
  wire  _T_19; // @[ALU.scala 70:41:freechips.rocketchip.system.DefaultRV32Config.fir@223161.4]
  wire [4:0] shamt; // @[ALU.scala 74:28:freechips.rocketchip.system.DefaultRV32Config.fir@223164.4]
  wire  _T_21; // @[ALU.scala 82:24:freechips.rocketchip.system.DefaultRV32Config.fir@223165.4]
  wire  _T_22; // @[ALU.scala 82:44:freechips.rocketchip.system.DefaultRV32Config.fir@223166.4]
  wire  _T_23; // @[ALU.scala 82:35:freechips.rocketchip.system.DefaultRV32Config.fir@223167.4]
  wire [31:0] _T_27; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@223171.4]
  wire [31:0] _T_29; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@223173.4]
  wire [31:0] _T_31; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@223175.4]
  wire [31:0] _T_32; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@223176.4]
  wire [31:0] _GEN_1; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@223181.4]
  wire [31:0] _T_37; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@223181.4]
  wire [31:0] _T_39; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@223183.4]
  wire [31:0] _T_41; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@223185.4]
  wire [31:0] _T_42; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@223186.4]
  wire [31:0] _GEN_2; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@223191.4]
  wire [31:0] _T_47; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@223191.4]
  wire [31:0] _T_49; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@223193.4]
  wire [31:0] _T_51; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@223195.4]
  wire [31:0] _T_52; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@223196.4]
  wire [31:0] _GEN_3; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@223201.4]
  wire [31:0] _T_57; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@223201.4]
  wire [31:0] _T_59; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@223203.4]
  wire [31:0] _T_61; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@223205.4]
  wire [31:0] _T_62; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@223206.4]
  wire [31:0] _GEN_4; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@223211.4]
  wire [31:0] _T_67; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@223211.4]
  wire [31:0] _T_69; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@223213.4]
  wire [31:0] _T_71; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@223215.4]
  wire [31:0] _T_72; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@223216.4]
  wire [31:0] shin; // @[ALU.scala 82:17:freechips.rocketchip.system.DefaultRV32Config.fir@223217.4]
  wire  _T_75; // @[ALU.scala 83:35:freechips.rocketchip.system.DefaultRV32Config.fir@223220.4]
  wire [32:0] _T_77; // @[ALU.scala 83:57:freechips.rocketchip.system.DefaultRV32Config.fir@223222.4]
  wire [32:0] _T_78; // @[ALU.scala 83:64:freechips.rocketchip.system.DefaultRV32Config.fir@223223.4]
  wire [31:0] shout_r; // @[ALU.scala 83:73:freechips.rocketchip.system.DefaultRV32Config.fir@223224.4]
  wire [31:0] _T_82; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@223228.4]
  wire [31:0] _T_84; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@223230.4]
  wire [31:0] _T_86; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@223232.4]
  wire [31:0] _T_87; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@223233.4]
  wire [31:0] _GEN_5; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@223238.4]
  wire [31:0] _T_92; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@223238.4]
  wire [31:0] _T_94; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@223240.4]
  wire [31:0] _T_96; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@223242.4]
  wire [31:0] _T_97; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@223243.4]
  wire [31:0] _GEN_6; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@223248.4]
  wire [31:0] _T_102; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@223248.4]
  wire [31:0] _T_104; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@223250.4]
  wire [31:0] _T_106; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@223252.4]
  wire [31:0] _T_107; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@223253.4]
  wire [31:0] _GEN_7; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@223258.4]
  wire [31:0] _T_112; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@223258.4]
  wire [31:0] _T_114; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@223260.4]
  wire [31:0] _T_116; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@223262.4]
  wire [31:0] _T_117; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@223263.4]
  wire [31:0] _GEN_8; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@223268.4]
  wire [31:0] _T_122; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@223268.4]
  wire [31:0] _T_124; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@223270.4]
  wire [31:0] _T_126; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@223272.4]
  wire [31:0] shout_l; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@223273.4]
  wire [31:0] _T_130; // @[ALU.scala 85:18:freechips.rocketchip.system.DefaultRV32Config.fir@223277.4]
  wire  _T_131; // @[ALU.scala 86:25:freechips.rocketchip.system.DefaultRV32Config.fir@223278.4]
  wire [31:0] _T_132; // @[ALU.scala 86:18:freechips.rocketchip.system.DefaultRV32Config.fir@223279.4]
  wire [31:0] shout; // @[ALU.scala 85:74:freechips.rocketchip.system.DefaultRV32Config.fir@223280.4]
  wire  _T_133; // @[ALU.scala 89:25:freechips.rocketchip.system.DefaultRV32Config.fir@223281.4]
  wire  _T_134; // @[ALU.scala 89:45:freechips.rocketchip.system.DefaultRV32Config.fir@223282.4]
  wire  _T_135; // @[ALU.scala 89:36:freechips.rocketchip.system.DefaultRV32Config.fir@223283.4]
  wire [31:0] _T_136; // @[ALU.scala 89:18:freechips.rocketchip.system.DefaultRV32Config.fir@223284.4]
  wire  _T_138; // @[ALU.scala 90:44:freechips.rocketchip.system.DefaultRV32Config.fir@223286.4]
  wire  _T_139; // @[ALU.scala 90:35:freechips.rocketchip.system.DefaultRV32Config.fir@223287.4]
  wire [31:0] _T_140; // @[ALU.scala 90:63:freechips.rocketchip.system.DefaultRV32Config.fir@223288.4]
  wire [31:0] _T_141; // @[ALU.scala 90:18:freechips.rocketchip.system.DefaultRV32Config.fir@223289.4]
  wire [31:0] logic_; // @[ALU.scala 89:78:freechips.rocketchip.system.DefaultRV32Config.fir@223290.4]
  wire  _T_142; // @[ALU.scala 41:30:freechips.rocketchip.system.DefaultRV32Config.fir@223291.4]
  wire  _T_143; // @[ALU.scala 91:35:freechips.rocketchip.system.DefaultRV32Config.fir@223292.4]
  wire [31:0] _GEN_9; // @[ALU.scala 91:43:freechips.rocketchip.system.DefaultRV32Config.fir@223293.4]
  wire [31:0] _T_144; // @[ALU.scala 91:43:freechips.rocketchip.system.DefaultRV32Config.fir@223293.4]
  wire [31:0] shift_logic; // @[ALU.scala 91:51:freechips.rocketchip.system.DefaultRV32Config.fir@223294.4]
  wire  _T_145; // @[ALU.scala 92:23:freechips.rocketchip.system.DefaultRV32Config.fir@223295.4]
  wire  _T_146; // @[ALU.scala 92:43:freechips.rocketchip.system.DefaultRV32Config.fir@223296.4]
  wire  _T_147; // @[ALU.scala 92:34:freechips.rocketchip.system.DefaultRV32Config.fir@223297.4]
  assign _T_1 = ~io_in2; // @[ALU.scala 62:35:freechips.rocketchip.system.DefaultRV32Config.fir@223139.4]
  assign in2_inv = io_fn[3] ? _T_1 : io_in2; // @[ALU.scala 62:20:freechips.rocketchip.system.DefaultRV32Config.fir@223140.4]
  assign in1_xor_in2 = io_in1 ^ in2_inv; // @[ALU.scala 63:28:freechips.rocketchip.system.DefaultRV32Config.fir@223141.4]
  assign _T_3 = io_in1 + in2_inv; // @[ALU.scala 64:26:freechips.rocketchip.system.DefaultRV32Config.fir@223143.4]
  assign _GEN_0 = {{31'd0}, io_fn[3]}; // @[ALU.scala 64:36:freechips.rocketchip.system.DefaultRV32Config.fir@223145.4]
  assign _T_9 = io_in1[31] == io_in2[31]; // @[ALU.scala 68:24:freechips.rocketchip.system.DefaultRV32Config.fir@223150.4]
  assign _T_14 = io_fn[1] ? io_in2[31] : io_in1[31]; // @[ALU.scala 69:8:freechips.rocketchip.system.DefaultRV32Config.fir@223155.4]
  assign slt = _T_9 ? io_adder_out[31] : _T_14; // @[ALU.scala 68:8:freechips.rocketchip.system.DefaultRV32Config.fir@223156.4]
  assign _T_17 = ~io_fn[3]; // @[ALU.scala 44:26:freechips.rocketchip.system.DefaultRV32Config.fir@223159.4]
  assign _T_18 = in1_xor_in2 == 32'h0; // @[ALU.scala 70:68:freechips.rocketchip.system.DefaultRV32Config.fir@223160.4]
  assign _T_19 = _T_17 ? _T_18 : slt; // @[ALU.scala 70:41:freechips.rocketchip.system.DefaultRV32Config.fir@223161.4]
  assign shamt = io_in2[4:0]; // @[ALU.scala 74:28:freechips.rocketchip.system.DefaultRV32Config.fir@223164.4]
  assign _T_21 = io_fn == 4'h5; // @[ALU.scala 82:24:freechips.rocketchip.system.DefaultRV32Config.fir@223165.4]
  assign _T_22 = io_fn == 4'hb; // @[ALU.scala 82:44:freechips.rocketchip.system.DefaultRV32Config.fir@223166.4]
  assign _T_23 = _T_21 | _T_22; // @[ALU.scala 82:35:freechips.rocketchip.system.DefaultRV32Config.fir@223167.4]
  assign _T_27 = {{16'd0}, io_in1[31:16]}; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@223171.4]
  assign _T_29 = {io_in1[15:0], 16'h0}; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@223173.4]
  assign _T_31 = _T_29 & 32'hffff0000; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@223175.4]
  assign _T_32 = _T_27 | _T_31; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@223176.4]
  assign _GEN_1 = {{8'd0}, _T_32[31:8]}; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@223181.4]
  assign _T_37 = _GEN_1 & 32'hff00ff; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@223181.4]
  assign _T_39 = {_T_32[23:0], 8'h0}; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@223183.4]
  assign _T_41 = _T_39 & 32'hff00ff00; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@223185.4]
  assign _T_42 = _T_37 | _T_41; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@223186.4]
  assign _GEN_2 = {{4'd0}, _T_42[31:4]}; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@223191.4]
  assign _T_47 = _GEN_2 & 32'hf0f0f0f; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@223191.4]
  assign _T_49 = {_T_42[27:0], 4'h0}; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@223193.4]
  assign _T_51 = _T_49 & 32'hf0f0f0f0; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@223195.4]
  assign _T_52 = _T_47 | _T_51; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@223196.4]
  assign _GEN_3 = {{2'd0}, _T_52[31:2]}; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@223201.4]
  assign _T_57 = _GEN_3 & 32'h33333333; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@223201.4]
  assign _T_59 = {_T_52[29:0], 2'h0}; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@223203.4]
  assign _T_61 = _T_59 & 32'hcccccccc; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@223205.4]
  assign _T_62 = _T_57 | _T_61; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@223206.4]
  assign _GEN_4 = {{1'd0}, _T_62[31:1]}; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@223211.4]
  assign _T_67 = _GEN_4 & 32'h55555555; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@223211.4]
  assign _T_69 = {_T_62[30:0], 1'h0}; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@223213.4]
  assign _T_71 = _T_69 & 32'haaaaaaaa; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@223215.4]
  assign _T_72 = _T_67 | _T_71; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@223216.4]
  assign shin = _T_23 ? io_in1 : _T_72; // @[ALU.scala 82:17:freechips.rocketchip.system.DefaultRV32Config.fir@223217.4]
  assign _T_75 = io_fn[3] & shin[31]; // @[ALU.scala 83:35:freechips.rocketchip.system.DefaultRV32Config.fir@223220.4]
  assign _T_77 = {_T_75,shin}; // @[ALU.scala 83:57:freechips.rocketchip.system.DefaultRV32Config.fir@223222.4]
  assign _T_78 = $signed(_T_77) >>> shamt; // @[ALU.scala 83:64:freechips.rocketchip.system.DefaultRV32Config.fir@223223.4]
  assign shout_r = _T_78[31:0]; // @[ALU.scala 83:73:freechips.rocketchip.system.DefaultRV32Config.fir@223224.4]
  assign _T_82 = {{16'd0}, shout_r[31:16]}; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@223228.4]
  assign _T_84 = {shout_r[15:0], 16'h0}; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@223230.4]
  assign _T_86 = _T_84 & 32'hffff0000; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@223232.4]
  assign _T_87 = _T_82 | _T_86; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@223233.4]
  assign _GEN_5 = {{8'd0}, _T_87[31:8]}; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@223238.4]
  assign _T_92 = _GEN_5 & 32'hff00ff; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@223238.4]
  assign _T_94 = {_T_87[23:0], 8'h0}; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@223240.4]
  assign _T_96 = _T_94 & 32'hff00ff00; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@223242.4]
  assign _T_97 = _T_92 | _T_96; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@223243.4]
  assign _GEN_6 = {{4'd0}, _T_97[31:4]}; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@223248.4]
  assign _T_102 = _GEN_6 & 32'hf0f0f0f; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@223248.4]
  assign _T_104 = {_T_97[27:0], 4'h0}; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@223250.4]
  assign _T_106 = _T_104 & 32'hf0f0f0f0; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@223252.4]
  assign _T_107 = _T_102 | _T_106; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@223253.4]
  assign _GEN_7 = {{2'd0}, _T_107[31:2]}; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@223258.4]
  assign _T_112 = _GEN_7 & 32'h33333333; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@223258.4]
  assign _T_114 = {_T_107[29:0], 2'h0}; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@223260.4]
  assign _T_116 = _T_114 & 32'hcccccccc; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@223262.4]
  assign _T_117 = _T_112 | _T_116; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@223263.4]
  assign _GEN_8 = {{1'd0}, _T_117[31:1]}; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@223268.4]
  assign _T_122 = _GEN_8 & 32'h55555555; // @[Bitwise.scala 103:31:freechips.rocketchip.system.DefaultRV32Config.fir@223268.4]
  assign _T_124 = {_T_117[30:0], 1'h0}; // @[Bitwise.scala 103:65:freechips.rocketchip.system.DefaultRV32Config.fir@223270.4]
  assign _T_126 = _T_124 & 32'haaaaaaaa; // @[Bitwise.scala 103:75:freechips.rocketchip.system.DefaultRV32Config.fir@223272.4]
  assign shout_l = _T_122 | _T_126; // @[Bitwise.scala 103:39:freechips.rocketchip.system.DefaultRV32Config.fir@223273.4]
  assign _T_130 = _T_23 ? shout_r : 32'h0; // @[ALU.scala 85:18:freechips.rocketchip.system.DefaultRV32Config.fir@223277.4]
  assign _T_131 = io_fn == 4'h1; // @[ALU.scala 86:25:freechips.rocketchip.system.DefaultRV32Config.fir@223278.4]
  assign _T_132 = _T_131 ? shout_l : 32'h0; // @[ALU.scala 86:18:freechips.rocketchip.system.DefaultRV32Config.fir@223279.4]
  assign shout = _T_130 | _T_132; // @[ALU.scala 85:74:freechips.rocketchip.system.DefaultRV32Config.fir@223280.4]
  assign _T_133 = io_fn == 4'h4; // @[ALU.scala 89:25:freechips.rocketchip.system.DefaultRV32Config.fir@223281.4]
  assign _T_134 = io_fn == 4'h6; // @[ALU.scala 89:45:freechips.rocketchip.system.DefaultRV32Config.fir@223282.4]
  assign _T_135 = _T_133 | _T_134; // @[ALU.scala 89:36:freechips.rocketchip.system.DefaultRV32Config.fir@223283.4]
  assign _T_136 = _T_135 ? in1_xor_in2 : 32'h0; // @[ALU.scala 89:18:freechips.rocketchip.system.DefaultRV32Config.fir@223284.4]
  assign _T_138 = io_fn == 4'h7; // @[ALU.scala 90:44:freechips.rocketchip.system.DefaultRV32Config.fir@223286.4]
  assign _T_139 = _T_134 | _T_138; // @[ALU.scala 90:35:freechips.rocketchip.system.DefaultRV32Config.fir@223287.4]
  assign _T_140 = io_in1 & io_in2; // @[ALU.scala 90:63:freechips.rocketchip.system.DefaultRV32Config.fir@223288.4]
  assign _T_141 = _T_139 ? _T_140 : 32'h0; // @[ALU.scala 90:18:freechips.rocketchip.system.DefaultRV32Config.fir@223289.4]
  assign logic_ = _T_136 | _T_141; // @[ALU.scala 89:78:freechips.rocketchip.system.DefaultRV32Config.fir@223290.4]
  assign _T_142 = io_fn >= 4'hc; // @[ALU.scala 41:30:freechips.rocketchip.system.DefaultRV32Config.fir@223291.4]
  assign _T_143 = _T_142 & slt; // @[ALU.scala 91:35:freechips.rocketchip.system.DefaultRV32Config.fir@223292.4]
  assign _GEN_9 = {{31'd0}, _T_143}; // @[ALU.scala 91:43:freechips.rocketchip.system.DefaultRV32Config.fir@223293.4]
  assign _T_144 = _GEN_9 | logic_; // @[ALU.scala 91:43:freechips.rocketchip.system.DefaultRV32Config.fir@223293.4]
  assign shift_logic = _T_144 | shout; // @[ALU.scala 91:51:freechips.rocketchip.system.DefaultRV32Config.fir@223294.4]
  assign _T_145 = io_fn == 4'h0; // @[ALU.scala 92:23:freechips.rocketchip.system.DefaultRV32Config.fir@223295.4]
  assign _T_146 = io_fn == 4'ha; // @[ALU.scala 92:43:freechips.rocketchip.system.DefaultRV32Config.fir@223296.4]
  assign _T_147 = _T_145 | _T_146; // @[ALU.scala 92:34:freechips.rocketchip.system.DefaultRV32Config.fir@223297.4]
  assign io_out = _T_147 ? io_adder_out : shift_logic; // @[ALU.scala 94:10:freechips.rocketchip.system.DefaultRV32Config.fir@223299.4]
  assign io_adder_out = _T_3 + _GEN_0; // @[ALU.scala 64:16:freechips.rocketchip.system.DefaultRV32Config.fir@223147.4]
  assign io_cmp_out = io_fn[0] ^ _T_19; // @[ALU.scala 70:14:freechips.rocketchip.system.DefaultRV32Config.fir@223163.4]
endmodule
