module TLMonitor_48( // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207509.2]
  input         clock, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207510.4]
  input         reset, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207511.4]
  input         io_in_a_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207512.4]
  input         io_in_a_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207512.4]
  input  [2:0]  io_in_a_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207512.4]
  input  [2:0]  io_in_a_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207512.4]
  input  [3:0]  io_in_a_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207512.4]
  input  [1:0]  io_in_a_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207512.4]
  input  [31:0] io_in_a_bits_address, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207512.4]
  input  [3:0]  io_in_a_bits_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207512.4]
  input         io_in_a_bits_corrupt, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207512.4]
  input         io_in_b_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207512.4]
  input         io_in_b_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207512.4]
  input  [2:0]  io_in_b_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207512.4]
  input  [1:0]  io_in_b_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207512.4]
  input  [3:0]  io_in_b_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207512.4]
  input  [1:0]  io_in_b_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207512.4]
  input  [31:0] io_in_b_bits_address, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207512.4]
  input  [3:0]  io_in_b_bits_mask, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207512.4]
  input         io_in_b_bits_corrupt, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207512.4]
  input         io_in_c_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207512.4]
  input         io_in_c_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207512.4]
  input  [2:0]  io_in_c_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207512.4]
  input  [2:0]  io_in_c_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207512.4]
  input  [3:0]  io_in_c_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207512.4]
  input  [1:0]  io_in_c_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207512.4]
  input  [31:0] io_in_c_bits_address, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207512.4]
  input         io_in_d_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207512.4]
  input         io_in_d_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207512.4]
  input  [2:0]  io_in_d_bits_opcode, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207512.4]
  input  [1:0]  io_in_d_bits_param, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207512.4]
  input  [3:0]  io_in_d_bits_size, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207512.4]
  input  [1:0]  io_in_d_bits_source, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207512.4]
  input  [1:0]  io_in_d_bits_sink, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207512.4]
  input         io_in_d_bits_denied, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207512.4]
  input         io_in_d_bits_corrupt, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207512.4]
  input         io_in_e_ready, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207512.4]
  input         io_in_e_valid, // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207512.4]
  input  [1:0]  io_in_e_bits_sink // @[:freechips.rocketchip.system.DefaultRV32Config.fir@207512.4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11:freechips.rocketchip.system.DefaultRV32Config.fir@210375.4]
  wire  _T_4; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@207523.6]
  wire  _T_5; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@207524.6]
  wire  _T_6; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@207525.6]
  wire  _T_8; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@207531.6]
  wire  _T_9; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@207532.6]
  wire [26:0] _T_11; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@207534.6]
  wire [11:0] _T_13; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@207536.6]
  wire [31:0] _GEN_71; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@207537.6]
  wire [31:0] _T_14; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@207537.6]
  wire  _T_15; // @[Edges.scala 22:24:freechips.rocketchip.system.DefaultRV32Config.fir@207538.6]
  wire [1:0] _T_18; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@207541.6]
  wire [1:0] _T_20; // @[Misc.scala 201:81:freechips.rocketchip.system.DefaultRV32Config.fir@207543.6]
  wire  _T_21; // @[Misc.scala 205:21:freechips.rocketchip.system.DefaultRV32Config.fir@207544.6]
  wire  _T_24; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@207547.6]
  wire  _T_26; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@207549.6]
  wire  _T_27; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@207550.6]
  wire  _T_29; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@207552.6]
  wire  _T_30; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@207553.6]
  wire  _T_33; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@207556.6]
  wire  _T_34; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@207557.6]
  wire  _T_35; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@207558.6]
  wire  _T_36; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@207559.6]
  wire  _T_37; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@207560.6]
  wire  _T_38; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@207561.6]
  wire  _T_39; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@207562.6]
  wire  _T_40; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@207563.6]
  wire  _T_41; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@207564.6]
  wire  _T_42; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@207565.6]
  wire  _T_43; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@207566.6]
  wire  _T_44; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@207567.6]
  wire  _T_45; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@207568.6]
  wire [3:0] _T_48; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@207571.6]
  wire [32:0] _T_52; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@207575.6]
  wire  _T_78; // @[Monitor.scala 79:25:freechips.rocketchip.system.DefaultRV32Config.fir@207605.6]
  wire [32:0] _T_83; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@207611.8]
  wire  _T_84; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@207612.8]
  wire [31:0] _T_85; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@207613.8]
  wire [32:0] _T_86; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@207614.8]
  wire [32:0] _T_88; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@207616.8]
  wire  _T_89; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@207617.8]
  wire [31:0] _T_90; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@207618.8]
  wire [32:0] _T_91; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@207619.8]
  wire [32:0] _T_93; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@207621.8]
  wire  _T_94; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@207622.8]
  wire [31:0] _T_95; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@207623.8]
  wire [32:0] _T_96; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@207624.8]
  wire [32:0] _T_98; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@207626.8]
  wire  _T_99; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@207627.8]
  wire [31:0] _T_100; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@207628.8]
  wire [32:0] _T_101; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@207629.8]
  wire [32:0] _T_103; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@207631.8]
  wire  _T_104; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@207632.8]
  wire [31:0] _T_105; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@207633.8]
  wire [32:0] _T_106; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@207634.8]
  wire [32:0] _T_108; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@207636.8]
  wire  _T_109; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@207637.8]
  wire  _T_110; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@207638.8]
  wire  _T_117; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@207645.8]
  wire [31:0] _T_120; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@207648.8]
  wire [32:0] _T_121; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@207649.8]
  wire [32:0] _T_123; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@207651.8]
  wire  _T_124; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@207652.8]
  wire  _T_125; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@207653.8]
  wire  _T_129; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207657.8]
  wire  _T_130; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207658.8]
  wire  _T_135; // @[Parameters.scala 92:48:freechips.rocketchip.system.DefaultRV32Config.fir@207671.8]
  wire  _T_136; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@207672.8]
  wire  _T_143; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207680.8]
  wire  _T_144; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207681.8]
  wire  _T_146; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207687.8]
  wire  _T_147; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207688.8]
  wire  _T_150; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207695.8]
  wire  _T_151; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207696.8]
  wire  _T_153; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207702.8]
  wire  _T_154; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207703.8]
  wire  _T_155; // @[Bundles.scala 110:27:freechips.rocketchip.system.DefaultRV32Config.fir@207708.8]
  wire  _T_157; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207710.8]
  wire  _T_158; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207711.8]
  wire [3:0] _T_159; // @[Monitor.scala 86:18:freechips.rocketchip.system.DefaultRV32Config.fir@207716.8]
  wire  _T_160; // @[Monitor.scala 86:31:freechips.rocketchip.system.DefaultRV32Config.fir@207717.8]
  wire  _T_162; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207719.8]
  wire  _T_163; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207720.8]
  wire  _T_164; // @[Monitor.scala 87:18:freechips.rocketchip.system.DefaultRV32Config.fir@207725.8]
  wire  _T_166; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207727.8]
  wire  _T_167; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207728.8]
  wire  _T_168; // @[Monitor.scala 90:25:freechips.rocketchip.system.DefaultRV32Config.fir@207734.6]
  wire  _T_249; // @[Monitor.scala 97:31:freechips.rocketchip.system.DefaultRV32Config.fir@207845.8]
  wire  _T_251; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207847.8]
  wire  _T_252; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207848.8]
  wire  _T_262; // @[Monitor.scala 102:25:freechips.rocketchip.system.DefaultRV32Config.fir@207871.6]
  wire  _T_264; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@207874.8]
  wire  _T_272; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@207882.8]
  wire  _T_307; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@207917.8]
  wire  _T_308; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@207918.8]
  wire  _T_309; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@207919.8]
  wire  _T_310; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@207920.8]
  wire  _T_311; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@207921.8]
  wire  _T_312; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@207922.8]
  wire  _T_314; // @[Parameters.scala 553:30:freechips.rocketchip.system.DefaultRV32Config.fir@207924.8]
  wire  _T_316; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207926.8]
  wire  _T_317; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207927.8]
  wire  _T_324; // @[Monitor.scala 106:31:freechips.rocketchip.system.DefaultRV32Config.fir@207946.8]
  wire  _T_326; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207948.8]
  wire  _T_327; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207949.8]
  wire  _T_328; // @[Monitor.scala 107:30:freechips.rocketchip.system.DefaultRV32Config.fir@207954.8]
  wire  _T_330; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207956.8]
  wire  _T_331; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207957.8]
  wire  _T_336; // @[Monitor.scala 111:25:freechips.rocketchip.system.DefaultRV32Config.fir@207971.6]
  wire  _T_371; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@208007.8]
  wire  _T_372; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@208008.8]
  wire  _T_373; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@208009.8]
  wire  _T_374; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@208010.8]
  wire  _T_383; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@208019.8]
  wire  _T_391; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@208027.8]
  wire  _T_393; // @[Parameters.scala 553:30:freechips.rocketchip.system.DefaultRV32Config.fir@208029.8]
  wire  _T_395; // @[Parameters.scala 553:30:freechips.rocketchip.system.DefaultRV32Config.fir@208031.8]
  wire  _T_397; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208033.8]
  wire  _T_398; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208034.8]
  wire  _T_413; // @[Monitor.scala 119:25:freechips.rocketchip.system.DefaultRV32Config.fir@208070.6]
  wire [3:0] _T_486; // @[Monitor.scala 124:33:freechips.rocketchip.system.DefaultRV32Config.fir@208160.8]
  wire [3:0] _T_487; // @[Monitor.scala 124:31:freechips.rocketchip.system.DefaultRV32Config.fir@208161.8]
  wire  _T_488; // @[Monitor.scala 124:40:freechips.rocketchip.system.DefaultRV32Config.fir@208162.8]
  wire  _T_490; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208164.8]
  wire  _T_491; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208165.8]
  wire  _T_492; // @[Monitor.scala 127:25:freechips.rocketchip.system.DefaultRV32Config.fir@208171.6]
  wire  _T_494; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@208174.8]
  wire  _T_518; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@208198.8]
  wire  _T_519; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@208199.8]
  wire  _T_520; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@208200.8]
  wire  _T_543; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208223.8]
  wire  _T_544; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208224.8]
  wire  _T_551; // @[Bundles.scala 140:33:freechips.rocketchip.system.DefaultRV32Config.fir@208243.8]
  wire  _T_553; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208245.8]
  wire  _T_554; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208246.8]
  wire  _T_559; // @[Monitor.scala 135:25:freechips.rocketchip.system.DefaultRV32Config.fir@208260.6]
  wire  _T_618; // @[Bundles.scala 147:30:freechips.rocketchip.system.DefaultRV32Config.fir@208332.8]
  wire  _T_620; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208334.8]
  wire  _T_621; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208335.8]
  wire  _T_626; // @[Monitor.scala 143:25:freechips.rocketchip.system.DefaultRV32Config.fir@208349.6]
  wire  _T_677; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208401.8]
  wire  _T_678; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208402.8]
  wire  _T_685; // @[Bundles.scala 160:28:freechips.rocketchip.system.DefaultRV32Config.fir@208421.8]
  wire  _T_687; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208423.8]
  wire  _T_688; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208424.8]
  wire  _T_697; // @[Bundles.scala 44:24:freechips.rocketchip.system.DefaultRV32Config.fir@208448.6]
  wire  _T_699; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208450.6]
  wire  _T_700; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208451.6]
  wire  _T_701; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@208456.6]
  wire  _T_702; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@208457.6]
  wire  _T_703; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@208458.6]
  wire  _T_705; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@208464.6]
  wire  _T_706; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@208465.6]
  wire  _T_708; // @[Monitor.scala 307:25:freechips.rocketchip.system.DefaultRV32Config.fir@208467.6]
  wire  _T_710; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208470.8]
  wire  _T_711; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208471.8]
  wire  _T_712; // @[Monitor.scala 309:27:freechips.rocketchip.system.DefaultRV32Config.fir@208476.8]
  wire  _T_714; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208478.8]
  wire  _T_715; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208479.8]
  wire  _T_716; // @[Monitor.scala 310:28:freechips.rocketchip.system.DefaultRV32Config.fir@208484.8]
  wire  _T_718; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208486.8]
  wire  _T_719; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208487.8]
  wire  _T_720; // @[Monitor.scala 311:15:freechips.rocketchip.system.DefaultRV32Config.fir@208492.8]
  wire  _T_722; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208494.8]
  wire  _T_723; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208495.8]
  wire  _T_724; // @[Monitor.scala 312:15:freechips.rocketchip.system.DefaultRV32Config.fir@208500.8]
  wire  _T_726; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208502.8]
  wire  _T_727; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208503.8]
  wire  _T_728; // @[Monitor.scala 315:25:freechips.rocketchip.system.DefaultRV32Config.fir@208509.6]
  wire  _T_739; // @[Bundles.scala 104:26:freechips.rocketchip.system.DefaultRV32Config.fir@208533.8]
  wire  _T_741; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208535.8]
  wire  _T_742; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208536.8]
  wire  _T_743; // @[Monitor.scala 320:28:freechips.rocketchip.system.DefaultRV32Config.fir@208541.8]
  wire  _T_745; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208543.8]
  wire  _T_746; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208544.8]
  wire  _T_756; // @[Monitor.scala 325:25:freechips.rocketchip.system.DefaultRV32Config.fir@208567.6]
  wire  _T_776; // @[Monitor.scala 331:30:freechips.rocketchip.system.DefaultRV32Config.fir@208608.8]
  wire  _T_778; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208610.8]
  wire  _T_779; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208611.8]
  wire  _T_785; // @[Monitor.scala 335:25:freechips.rocketchip.system.DefaultRV32Config.fir@208626.6]
  wire  _T_802; // @[Monitor.scala 343:25:freechips.rocketchip.system.DefaultRV32Config.fir@208661.6]
  wire  _T_820; // @[Monitor.scala 351:25:freechips.rocketchip.system.DefaultRV32Config.fir@208697.6]
  wire  _T_837; // @[Bundles.scala 42:24:freechips.rocketchip.system.DefaultRV32Config.fir@208734.6]
  wire  _T_839; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208736.6]
  wire  _T_840; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208737.6]
  wire  _T_841; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@208742.6]
  wire [32:0] _T_844; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208745.6]
  wire  _T_849; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@208750.6]
  wire  _T_857; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@208758.6]
  wire [31:0] _T_870; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@208775.6]
  wire [32:0] _T_871; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208776.6]
  wire [32:0] _T_873; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208778.6]
  wire  _T_874; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208779.6]
  wire [31:0] _T_875; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@208780.6]
  wire [32:0] _T_876; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208781.6]
  wire [32:0] _T_878; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208783.6]
  wire  _T_879; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208784.6]
  wire [31:0] _T_880; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@208785.6]
  wire [32:0] _T_881; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208786.6]
  wire [32:0] _T_883; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208788.6]
  wire  _T_884; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208789.6]
  wire [32:0] _T_888; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208793.6]
  wire  _T_889; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208794.6]
  wire [31:0] _T_890; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@208795.6]
  wire [32:0] _T_891; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208796.6]
  wire [32:0] _T_893; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208798.6]
  wire  _T_894; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208799.6]
  wire [31:0] _T_895; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@208800.6]
  wire [32:0] _T_896; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208801.6]
  wire [32:0] _T_898; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208803.6]
  wire  _T_899; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208804.6]
  wire [31:0] _T_900; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@208805.6]
  wire [32:0] _T_901; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208806.6]
  wire [32:0] _T_903; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208808.6]
  wire  _T_904; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208809.6]
  wire  _T_906; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@208819.6]
  wire  _T_907; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@208820.6]
  wire  _T_908; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@208821.6]
  wire  _T_909; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@208822.6]
  wire  _T_910; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@208823.6]
  wire  _T_911; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@208824.6]
  wire [26:0] _T_913; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@208826.6]
  wire [11:0] _T_915; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@208828.6]
  wire [31:0] _GEN_72; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@208829.6]
  wire [31:0] _T_916; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@208829.6]
  wire  _T_917; // @[Edges.scala 22:24:freechips.rocketchip.system.DefaultRV32Config.fir@208830.6]
  wire [1:0] _T_920; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@208833.6]
  wire [1:0] _T_922; // @[Misc.scala 201:81:freechips.rocketchip.system.DefaultRV32Config.fir@208835.6]
  wire  _T_923; // @[Misc.scala 205:21:freechips.rocketchip.system.DefaultRV32Config.fir@208836.6]
  wire  _T_926; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@208839.6]
  wire  _T_928; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@208841.6]
  wire  _T_929; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@208842.6]
  wire  _T_931; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@208844.6]
  wire  _T_932; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@208845.6]
  wire  _T_935; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@208848.6]
  wire  _T_936; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@208849.6]
  wire  _T_937; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@208850.6]
  wire  _T_938; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@208851.6]
  wire  _T_939; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@208852.6]
  wire  _T_940; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@208853.6]
  wire  _T_941; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@208854.6]
  wire  _T_942; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@208855.6]
  wire  _T_943; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@208856.6]
  wire  _T_944; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@208857.6]
  wire  _T_945; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@208858.6]
  wire  _T_946; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@208859.6]
  wire  _T_947; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@208860.6]
  wire [3:0] _T_950; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@208863.6]
  wire [1:0] _T_957; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@208874.6]
  wire [1:0] _GEN_73; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@208876.6]
  wire [1:0] _T_959; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@208876.6]
  wire  _T_961; // @[Monitor.scala 162:113:freechips.rocketchip.system.DefaultRV32Config.fir@208879.6]
  wire  _T_962; // @[Monitor.scala 164:25:freechips.rocketchip.system.DefaultRV32Config.fir@208880.6]
  wire  _T_967; // @[Parameters.scala 92:48:freechips.rocketchip.system.DefaultRV32Config.fir@208890.8]
  wire  _T_968; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@208891.8]
  wire  _T_975; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208899.8]
  wire  _T_976; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208900.8]
  wire  _T_978; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208906.8]
  wire  _T_979; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208907.8]
  wire  _T_981; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208913.8]
  wire  _T_982; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208914.8]
  wire  _T_984; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208920.8]
  wire  _T_985; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208921.8]
  wire  _T_986; // @[Bundles.scala 104:26:freechips.rocketchip.system.DefaultRV32Config.fir@208926.8]
  wire  _T_988; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208928.8]
  wire  _T_989; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208929.8]
  wire  _T_990; // @[Monitor.scala 170:30:freechips.rocketchip.system.DefaultRV32Config.fir@208934.8]
  wire  _T_992; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208936.8]
  wire  _T_993; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208937.8]
  wire  _T_994; // @[Monitor.scala 171:18:freechips.rocketchip.system.DefaultRV32Config.fir@208942.8]
  wire  _T_996; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208944.8]
  wire  _T_997; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208945.8]
  wire  _T_998; // @[Monitor.scala 174:25:freechips.rocketchip.system.DefaultRV32Config.fir@208951.6]
  wire  _T_1001; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208955.8]
  wire  _T_1011; // @[Monitor.scala 179:31:freechips.rocketchip.system.DefaultRV32Config.fir@208981.8]
  wire  _T_1013; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208983.8]
  wire  _T_1014; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208984.8]
  wire  _T_1023; // @[Monitor.scala 184:25:freechips.rocketchip.system.DefaultRV32Config.fir@209006.6]
  wire  _T_1044; // @[Monitor.scala 193:25:freechips.rocketchip.system.DefaultRV32Config.fir@209053.6]
  wire [3:0] _T_1061; // @[Monitor.scala 199:33:freechips.rocketchip.system.DefaultRV32Config.fir@209091.8]
  wire [3:0] _T_1062; // @[Monitor.scala 199:31:freechips.rocketchip.system.DefaultRV32Config.fir@209092.8]
  wire  _T_1063; // @[Monitor.scala 199:40:freechips.rocketchip.system.DefaultRV32Config.fir@209093.8]
  wire  _T_1065; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209095.8]
  wire  _T_1066; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209096.8]
  wire  _T_1067; // @[Monitor.scala 202:25:freechips.rocketchip.system.DefaultRV32Config.fir@209102.6]
  wire  _T_1088; // @[Monitor.scala 211:25:freechips.rocketchip.system.DefaultRV32Config.fir@209149.6]
  wire  _T_1109; // @[Monitor.scala 220:25:freechips.rocketchip.system.DefaultRV32Config.fir@209196.6]
  wire  _T_1134; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@209253.6]
  wire  _T_1135; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@209254.6]
  wire  _T_1136; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@209255.6]
  wire  _T_1138; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@209261.6]
  wire  _T_1139; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@209262.6]
  wire [26:0] _T_1141; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@209264.6]
  wire [11:0] _T_1143; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@209266.6]
  wire [31:0] _GEN_74; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@209267.6]
  wire [31:0] _T_1144; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@209267.6]
  wire  _T_1145; // @[Edges.scala 22:24:freechips.rocketchip.system.DefaultRV32Config.fir@209268.6]
  wire [31:0] _T_1146; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@209269.6]
  wire [32:0] _T_1147; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@209270.6]
  wire [32:0] _T_1149; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@209272.6]
  wire  _T_1150; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@209273.6]
  wire [31:0] _T_1151; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@209274.6]
  wire [32:0] _T_1152; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@209275.6]
  wire [32:0] _T_1154; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@209277.6]
  wire  _T_1155; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@209278.6]
  wire [31:0] _T_1156; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@209279.6]
  wire [32:0] _T_1157; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@209280.6]
  wire [32:0] _T_1159; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@209282.6]
  wire  _T_1160; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@209283.6]
  wire [32:0] _T_1162; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@209285.6]
  wire [32:0] _T_1164; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@209287.6]
  wire  _T_1165; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@209288.6]
  wire [31:0] _T_1166; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@209289.6]
  wire [32:0] _T_1167; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@209290.6]
  wire [32:0] _T_1169; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@209292.6]
  wire  _T_1170; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@209293.6]
  wire [31:0] _T_1171; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@209294.6]
  wire [32:0] _T_1172; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@209295.6]
  wire [32:0] _T_1174; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@209297.6]
  wire  _T_1175; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@209298.6]
  wire [31:0] _T_1176; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@209299.6]
  wire [32:0] _T_1177; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@209300.6]
  wire [32:0] _T_1179; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@209302.6]
  wire  _T_1180; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@209303.6]
  wire  _T_1182; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@209313.6]
  wire  _T_1183; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@209314.6]
  wire  _T_1184; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@209315.6]
  wire  _T_1185; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@209316.6]
  wire  _T_1186; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@209317.6]
  wire  _T_1187; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@209318.6]
  wire  _T_1217; // @[Monitor.scala 239:25:freechips.rocketchip.system.DefaultRV32Config.fir@209352.6]
  wire  _T_1219; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209355.8]
  wire  _T_1220; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209356.8]
  wire  _T_1222; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209362.8]
  wire  _T_1223; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209363.8]
  wire  _T_1224; // @[Monitor.scala 242:30:freechips.rocketchip.system.DefaultRV32Config.fir@209368.8]
  wire  _T_1226; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209370.8]
  wire  _T_1227; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209371.8]
  wire  _T_1229; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209377.8]
  wire  _T_1230; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209378.8]
  wire  _T_1231; // @[Bundles.scala 122:29:freechips.rocketchip.system.DefaultRV32Config.fir@209383.8]
  wire  _T_1233; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209385.8]
  wire  _T_1234; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209386.8]
  wire  _T_1239; // @[Monitor.scala 248:25:freechips.rocketchip.system.DefaultRV32Config.fir@209400.6]
  wire  _T_1257; // @[Monitor.scala 256:25:freechips.rocketchip.system.DefaultRV32Config.fir@209440.6]
  wire  _T_1296; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@209480.8]
  wire  _T_1304; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@209488.8]
  wire  _T_1308; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209492.8]
  wire  _T_1309; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209493.8]
  wire  _T_1314; // @[Parameters.scala 92:48:freechips.rocketchip.system.DefaultRV32Config.fir@209506.8]
  wire  _T_1315; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@209507.8]
  wire  _T_1322; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209515.8]
  wire  _T_1323; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209516.8]
  wire  _T_1334; // @[Bundles.scala 116:29:freechips.rocketchip.system.DefaultRV32Config.fir@209543.8]
  wire  _T_1336; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209545.8]
  wire  _T_1337; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209546.8]
  wire  _T_1342; // @[Monitor.scala 266:25:freechips.rocketchip.system.DefaultRV32Config.fir@209560.6]
  wire  _T_1423; // @[Monitor.scala 275:25:freechips.rocketchip.system.DefaultRV32Config.fir@209672.6]
  wire  _T_1433; // @[Monitor.scala 279:31:freechips.rocketchip.system.DefaultRV32Config.fir@209695.8]
  wire  _T_1435; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209697.8]
  wire  _T_1436; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209698.8]
  wire  _T_1441; // @[Monitor.scala 283:25:freechips.rocketchip.system.DefaultRV32Config.fir@209712.6]
  wire  _T_1455; // @[Monitor.scala 290:25:freechips.rocketchip.system.DefaultRV32Config.fir@209744.6]
  wire  _T_1477; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@209795.4]
  wire  _T_1484; // @[Edges.scala 93:28:freechips.rocketchip.system.DefaultRV32Config.fir@209802.4]
  reg [9:0] _T_1486; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@209804.4]
  wire [9:0] _T_1488; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@209806.4]
  wire  _T_1489; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@209807.4]
  reg [2:0] _T_1497; // @[Monitor.scala 381:22:freechips.rocketchip.system.DefaultRV32Config.fir@209818.4]
  reg [2:0] _T_1498; // @[Monitor.scala 382:22:freechips.rocketchip.system.DefaultRV32Config.fir@209819.4]
  reg [3:0] _T_1499; // @[Monitor.scala 383:22:freechips.rocketchip.system.DefaultRV32Config.fir@209820.4]
  reg [1:0] _T_1500; // @[Monitor.scala 384:22:freechips.rocketchip.system.DefaultRV32Config.fir@209821.4]
  reg [31:0] _T_1501; // @[Monitor.scala 385:22:freechips.rocketchip.system.DefaultRV32Config.fir@209822.4]
  wire  _T_1502; // @[Monitor.scala 386:22:freechips.rocketchip.system.DefaultRV32Config.fir@209823.4]
  wire  _T_1503; // @[Monitor.scala 386:19:freechips.rocketchip.system.DefaultRV32Config.fir@209824.4]
  wire  _T_1504; // @[Monitor.scala 387:32:freechips.rocketchip.system.DefaultRV32Config.fir@209826.6]
  wire  _T_1506; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209828.6]
  wire  _T_1507; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209829.6]
  wire  _T_1508; // @[Monitor.scala 388:32:freechips.rocketchip.system.DefaultRV32Config.fir@209834.6]
  wire  _T_1510; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209836.6]
  wire  _T_1511; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209837.6]
  wire  _T_1512; // @[Monitor.scala 389:32:freechips.rocketchip.system.DefaultRV32Config.fir@209842.6]
  wire  _T_1514; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209844.6]
  wire  _T_1515; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209845.6]
  wire  _T_1516; // @[Monitor.scala 390:32:freechips.rocketchip.system.DefaultRV32Config.fir@209850.6]
  wire  _T_1518; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209852.6]
  wire  _T_1519; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209853.6]
  wire  _T_1520; // @[Monitor.scala 391:32:freechips.rocketchip.system.DefaultRV32Config.fir@209858.6]
  wire  _T_1522; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209860.6]
  wire  _T_1523; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209861.6]
  wire  _T_1525; // @[Monitor.scala 393:20:freechips.rocketchip.system.DefaultRV32Config.fir@209868.4]
  wire  _T_1526; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@209876.4]
  wire [26:0] _T_1528; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@209878.4]
  wire [11:0] _T_1530; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@209880.4]
  reg [9:0] _T_1534; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@209884.4]
  wire [9:0] _T_1536; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@209886.4]
  wire  _T_1537; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@209887.4]
  reg [2:0] _T_1545; // @[Monitor.scala 532:22:freechips.rocketchip.system.DefaultRV32Config.fir@209898.4]
  reg [1:0] _T_1546; // @[Monitor.scala 533:22:freechips.rocketchip.system.DefaultRV32Config.fir@209899.4]
  reg [3:0] _T_1547; // @[Monitor.scala 534:22:freechips.rocketchip.system.DefaultRV32Config.fir@209900.4]
  reg [1:0] _T_1548; // @[Monitor.scala 535:22:freechips.rocketchip.system.DefaultRV32Config.fir@209901.4]
  reg [1:0] _T_1549; // @[Monitor.scala 536:22:freechips.rocketchip.system.DefaultRV32Config.fir@209902.4]
  reg  _T_1550; // @[Monitor.scala 537:22:freechips.rocketchip.system.DefaultRV32Config.fir@209903.4]
  wire  _T_1551; // @[Monitor.scala 538:22:freechips.rocketchip.system.DefaultRV32Config.fir@209904.4]
  wire  _T_1552; // @[Monitor.scala 538:19:freechips.rocketchip.system.DefaultRV32Config.fir@209905.4]
  wire  _T_1553; // @[Monitor.scala 539:29:freechips.rocketchip.system.DefaultRV32Config.fir@209907.6]
  wire  _T_1555; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209909.6]
  wire  _T_1556; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209910.6]
  wire  _T_1557; // @[Monitor.scala 540:29:freechips.rocketchip.system.DefaultRV32Config.fir@209915.6]
  wire  _T_1559; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209917.6]
  wire  _T_1560; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209918.6]
  wire  _T_1561; // @[Monitor.scala 541:29:freechips.rocketchip.system.DefaultRV32Config.fir@209923.6]
  wire  _T_1563; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209925.6]
  wire  _T_1564; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209926.6]
  wire  _T_1565; // @[Monitor.scala 542:29:freechips.rocketchip.system.DefaultRV32Config.fir@209931.6]
  wire  _T_1567; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209933.6]
  wire  _T_1568; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209934.6]
  wire  _T_1569; // @[Monitor.scala 543:29:freechips.rocketchip.system.DefaultRV32Config.fir@209939.6]
  wire  _T_1571; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209941.6]
  wire  _T_1572; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209942.6]
  wire  _T_1573; // @[Monitor.scala 544:29:freechips.rocketchip.system.DefaultRV32Config.fir@209947.6]
  wire  _T_1575; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209949.6]
  wire  _T_1576; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209950.6]
  wire  _T_1578; // @[Monitor.scala 546:20:freechips.rocketchip.system.DefaultRV32Config.fir@209957.4]
  wire  _T_1579; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@209966.4]
  reg [9:0] _T_1588; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@209975.4]
  wire [9:0] _T_1590; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@209977.4]
  wire  _T_1591; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@209978.4]
  reg [2:0] _T_1599; // @[Monitor.scala 404:22:freechips.rocketchip.system.DefaultRV32Config.fir@209989.4]
  reg [1:0] _T_1600; // @[Monitor.scala 405:22:freechips.rocketchip.system.DefaultRV32Config.fir@209990.4]
  reg [3:0] _T_1601; // @[Monitor.scala 406:22:freechips.rocketchip.system.DefaultRV32Config.fir@209991.4]
  reg [1:0] _T_1602; // @[Monitor.scala 407:22:freechips.rocketchip.system.DefaultRV32Config.fir@209992.4]
  reg [31:0] _T_1603; // @[Monitor.scala 408:22:freechips.rocketchip.system.DefaultRV32Config.fir@209993.4]
  wire  _T_1604; // @[Monitor.scala 409:22:freechips.rocketchip.system.DefaultRV32Config.fir@209994.4]
  wire  _T_1605; // @[Monitor.scala 409:19:freechips.rocketchip.system.DefaultRV32Config.fir@209995.4]
  wire  _T_1606; // @[Monitor.scala 410:32:freechips.rocketchip.system.DefaultRV32Config.fir@209997.6]
  wire  _T_1608; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209999.6]
  wire  _T_1609; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210000.6]
  wire  _T_1610; // @[Monitor.scala 411:32:freechips.rocketchip.system.DefaultRV32Config.fir@210005.6]
  wire  _T_1612; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210007.6]
  wire  _T_1613; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210008.6]
  wire  _T_1614; // @[Monitor.scala 412:32:freechips.rocketchip.system.DefaultRV32Config.fir@210013.6]
  wire  _T_1616; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210015.6]
  wire  _T_1617; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210016.6]
  wire  _T_1618; // @[Monitor.scala 413:32:freechips.rocketchip.system.DefaultRV32Config.fir@210021.6]
  wire  _T_1620; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210023.6]
  wire  _T_1621; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210024.6]
  wire  _T_1622; // @[Monitor.scala 414:32:freechips.rocketchip.system.DefaultRV32Config.fir@210029.6]
  wire  _T_1624; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210031.6]
  wire  _T_1625; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210032.6]
  wire  _T_1627; // @[Monitor.scala 416:20:freechips.rocketchip.system.DefaultRV32Config.fir@210039.4]
  wire  _T_1628; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@210047.4]
  reg [9:0] _T_1636; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@210055.4]
  wire [9:0] _T_1638; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@210057.4]
  wire  _T_1639; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@210058.4]
  reg [2:0] _T_1647; // @[Monitor.scala 509:22:freechips.rocketchip.system.DefaultRV32Config.fir@210069.4]
  reg [2:0] _T_1648; // @[Monitor.scala 510:22:freechips.rocketchip.system.DefaultRV32Config.fir@210070.4]
  reg [3:0] _T_1649; // @[Monitor.scala 511:22:freechips.rocketchip.system.DefaultRV32Config.fir@210071.4]
  reg [1:0] _T_1650; // @[Monitor.scala 512:22:freechips.rocketchip.system.DefaultRV32Config.fir@210072.4]
  reg [31:0] _T_1651; // @[Monitor.scala 513:22:freechips.rocketchip.system.DefaultRV32Config.fir@210073.4]
  wire  _T_1652; // @[Monitor.scala 514:22:freechips.rocketchip.system.DefaultRV32Config.fir@210074.4]
  wire  _T_1653; // @[Monitor.scala 514:19:freechips.rocketchip.system.DefaultRV32Config.fir@210075.4]
  wire  _T_1654; // @[Monitor.scala 515:32:freechips.rocketchip.system.DefaultRV32Config.fir@210077.6]
  wire  _T_1656; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210079.6]
  wire  _T_1657; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210080.6]
  wire  _T_1658; // @[Monitor.scala 516:32:freechips.rocketchip.system.DefaultRV32Config.fir@210085.6]
  wire  _T_1660; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210087.6]
  wire  _T_1661; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210088.6]
  wire  _T_1662; // @[Monitor.scala 517:32:freechips.rocketchip.system.DefaultRV32Config.fir@210093.6]
  wire  _T_1664; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210095.6]
  wire  _T_1665; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210096.6]
  wire  _T_1666; // @[Monitor.scala 518:32:freechips.rocketchip.system.DefaultRV32Config.fir@210101.6]
  wire  _T_1668; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210103.6]
  wire  _T_1669; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210104.6]
  wire  _T_1670; // @[Monitor.scala 519:32:freechips.rocketchip.system.DefaultRV32Config.fir@210109.6]
  wire  _T_1672; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210111.6]
  wire  _T_1673; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210112.6]
  wire  _T_1675; // @[Monitor.scala 521:20:freechips.rocketchip.system.DefaultRV32Config.fir@210119.4]
  reg [2:0] inflight; // @[Monitor.scala 608:27:freechips.rocketchip.system.DefaultRV32Config.fir@210127.4]
  reg [11:0] inflight_opcodes; // @[Monitor.scala 610:35:freechips.rocketchip.system.DefaultRV32Config.fir@210128.4]
  reg [23:0] inflight_sizes; // @[Monitor.scala 612:33:freechips.rocketchip.system.DefaultRV32Config.fir@210129.4]
  reg [9:0] _T_1685; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@210139.4]
  wire [9:0] _T_1687; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@210141.4]
  wire  a_first; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@210142.4]
  reg [9:0] _T_1703; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@210161.4]
  wire [9:0] _T_1705; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@210163.4]
  wire  d_first; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@210164.4]
  wire [3:0] _GEN_75; // @[Monitor.scala 629:69:freechips.rocketchip.system.DefaultRV32Config.fir@210183.4]
  wire [4:0] _T_1713; // @[Monitor.scala 629:69:freechips.rocketchip.system.DefaultRV32Config.fir@210183.4]
  wire [11:0] _T_1714; // @[Monitor.scala 629:44:freechips.rocketchip.system.DefaultRV32Config.fir@210184.4]
  wire [15:0] _T_1718; // @[Monitor.scala 606:57:freechips.rocketchip.system.DefaultRV32Config.fir@210188.4]
  wire [15:0] _GEN_76; // @[Monitor.scala 629:97:freechips.rocketchip.system.DefaultRV32Config.fir@210189.4]
  wire [15:0] _T_1719; // @[Monitor.scala 629:97:freechips.rocketchip.system.DefaultRV32Config.fir@210189.4]
  wire [15:0] _T_1720; // @[Monitor.scala 629:152:freechips.rocketchip.system.DefaultRV32Config.fir@210190.4]
  wire [4:0] _T_1721; // @[Monitor.scala 633:65:freechips.rocketchip.system.DefaultRV32Config.fir@210194.4]
  wire [23:0] _T_1722; // @[Monitor.scala 633:40:freechips.rocketchip.system.DefaultRV32Config.fir@210195.4]
  wire [15:0] _T_1726; // @[Monitor.scala 606:57:freechips.rocketchip.system.DefaultRV32Config.fir@210199.4]
  wire [23:0] _GEN_78; // @[Monitor.scala 633:91:freechips.rocketchip.system.DefaultRV32Config.fir@210200.4]
  wire [23:0] _T_1727; // @[Monitor.scala 633:91:freechips.rocketchip.system.DefaultRV32Config.fir@210200.4]
  wire [23:0] _T_1728; // @[Monitor.scala 633:144:freechips.rocketchip.system.DefaultRV32Config.fir@210201.4]
  wire  _T_1732; // @[Monitor.scala 643:27:freechips.rocketchip.system.DefaultRV32Config.fir@210226.4]
  wire [3:0] _T_1734; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@210229.6]
  wire [3:0] _T_1735; // @[Monitor.scala 645:53:freechips.rocketchip.system.DefaultRV32Config.fir@210231.6]
  wire [3:0] _T_1736; // @[Monitor.scala 645:61:freechips.rocketchip.system.DefaultRV32Config.fir@210232.6]
  wire [4:0] _T_1737; // @[Monitor.scala 646:49:freechips.rocketchip.system.DefaultRV32Config.fir@210234.6]
  wire [4:0] _T_1738; // @[Monitor.scala 646:57:freechips.rocketchip.system.DefaultRV32Config.fir@210235.6]
  wire [3:0] _GEN_80; // @[Monitor.scala 647:72:freechips.rocketchip.system.DefaultRV32Config.fir@210237.6]
  wire [4:0] _T_1739; // @[Monitor.scala 647:72:freechips.rocketchip.system.DefaultRV32Config.fir@210237.6]
  wire [3:0] a_opcodes_set_interm; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@210228.4]
  wire [34:0] _GEN_81; // @[Monitor.scala 647:47:freechips.rocketchip.system.DefaultRV32Config.fir@210238.6]
  wire [34:0] _T_1740; // @[Monitor.scala 647:47:freechips.rocketchip.system.DefaultRV32Config.fir@210238.6]
  wire [4:0] _T_1741; // @[Monitor.scala 648:68:freechips.rocketchip.system.DefaultRV32Config.fir@210240.6]
  wire [4:0] a_sizes_set_interm; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@210228.4]
  wire [35:0] _GEN_82; // @[Monitor.scala 648:43:freechips.rocketchip.system.DefaultRV32Config.fir@210241.6]
  wire [35:0] _T_1742; // @[Monitor.scala 648:43:freechips.rocketchip.system.DefaultRV32Config.fir@210241.6]
  wire [2:0] _T_1743; // @[Monitor.scala 649:26:freechips.rocketchip.system.DefaultRV32Config.fir@210243.6]
  wire  _T_1745; // @[Monitor.scala 649:17:freechips.rocketchip.system.DefaultRV32Config.fir@210245.6]
  wire  _T_1747; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210247.6]
  wire  _T_1748; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210248.6]
  wire [3:0] _GEN_27; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@210228.4]
  wire [34:0] _GEN_30; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@210228.4]
  wire [35:0] _GEN_31; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@210228.4]
  wire  _T_1751; // @[Monitor.scala 660:27:freechips.rocketchip.system.DefaultRV32Config.fir@210262.4]
  wire  _T_1753; // @[Monitor.scala 660:75:freechips.rocketchip.system.DefaultRV32Config.fir@210264.4]
  wire  _T_1754; // @[Monitor.scala 660:72:freechips.rocketchip.system.DefaultRV32Config.fir@210265.4]
  wire [3:0] _T_1755; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@210267.6]
  wire [46:0] _GEN_84; // @[Monitor.scala 662:76:freechips.rocketchip.system.DefaultRV32Config.fir@210274.6]
  wire [46:0] _T_1761; // @[Monitor.scala 662:76:freechips.rocketchip.system.DefaultRV32Config.fir@210274.6]
  wire [46:0] _GEN_85; // @[Monitor.scala 663:72:freechips.rocketchip.system.DefaultRV32Config.fir@210281.6]
  wire [46:0] _T_1767; // @[Monitor.scala 663:72:freechips.rocketchip.system.DefaultRV32Config.fir@210281.6]
  wire [3:0] _GEN_32; // @[Monitor.scala 660:91:freechips.rocketchip.system.DefaultRV32Config.fir@210266.4]
  wire [46:0] _GEN_33; // @[Monitor.scala 660:91:freechips.rocketchip.system.DefaultRV32Config.fir@210266.4]
  wire [46:0] _GEN_34; // @[Monitor.scala 660:91:freechips.rocketchip.system.DefaultRV32Config.fir@210266.4]
  wire  _T_1768; // @[Monitor.scala 665:26:freechips.rocketchip.system.DefaultRV32Config.fir@210284.4]
  wire  _T_1771; // @[Monitor.scala 665:71:freechips.rocketchip.system.DefaultRV32Config.fir@210287.4]
  wire [2:0] _T_1772; // @[Monitor.scala 666:25:freechips.rocketchip.system.DefaultRV32Config.fir@210289.6]
  wire  _T_1774; // @[Monitor.scala 666:93:freechips.rocketchip.system.DefaultRV32Config.fir@210291.6]
  wire  _T_1775; // @[Monitor.scala 666:68:freechips.rocketchip.system.DefaultRV32Config.fir@210292.6]
  wire  _T_1776; // @[Monitor.scala 666:142:freechips.rocketchip.system.DefaultRV32Config.fir@210293.6]
  wire  _T_1777; // @[Monitor.scala 666:119:freechips.rocketchip.system.DefaultRV32Config.fir@210294.6]
  wire  _T_1778; // @[Monitor.scala 666:166:freechips.rocketchip.system.DefaultRV32Config.fir@210295.6]
  wire  _T_1779; // @[Monitor.scala 666:49:freechips.rocketchip.system.DefaultRV32Config.fir@210296.6]
  wire  _T_1781; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210298.6]
  wire  _T_1782; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210299.6]
  wire [3:0] a_opcode_lookup; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@210181.4 :freechips.rocketchip.system.DefaultRV32Config.fir@210182.4 Monitor.scala 629:21:freechips.rocketchip.system.DefaultRV32Config.fir@210191.4]
  wire [2:0] _GEN_37; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@210305.6]
  wire [2:0] _GEN_38; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@210305.6]
  wire [2:0] _GEN_39; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@210305.6]
  wire [2:0] _GEN_40; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@210305.6]
  wire [2:0] _GEN_41; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@210305.6]
  wire [2:0] _GEN_42; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@210305.6]
  wire  _T_1784; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@210305.6]
  wire [2:0] _GEN_49; // @[Monitor.scala 667:96:freechips.rocketchip.system.DefaultRV32Config.fir@210307.6]
  wire [2:0] _GEN_50; // @[Monitor.scala 667:96:freechips.rocketchip.system.DefaultRV32Config.fir@210307.6]
  wire  _T_1786; // @[Monitor.scala 667:96:freechips.rocketchip.system.DefaultRV32Config.fir@210307.6]
  wire  _T_1787; // @[Monitor.scala 667:71:freechips.rocketchip.system.DefaultRV32Config.fir@210308.6]
  wire [2:0] _GEN_53; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@210309.6]
  wire [2:0] _GEN_54; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@210309.6]
  wire [2:0] _GEN_55; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@210309.6]
  wire [2:0] _GEN_56; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@210309.6]
  wire [2:0] _GEN_57; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@210309.6]
  wire [2:0] _GEN_58; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@210309.6]
  wire  _T_1788; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@210309.6]
  wire [2:0] _GEN_65; // @[Monitor.scala 668:124:freechips.rocketchip.system.DefaultRV32Config.fir@210310.6]
  wire [2:0] _GEN_66; // @[Monitor.scala 668:124:freechips.rocketchip.system.DefaultRV32Config.fir@210310.6]
  wire  _T_1789; // @[Monitor.scala 668:124:freechips.rocketchip.system.DefaultRV32Config.fir@210310.6]
  wire  _T_1790; // @[Monitor.scala 668:99:freechips.rocketchip.system.DefaultRV32Config.fir@210311.6]
  wire  _T_1791; // @[Monitor.scala 668:34:freechips.rocketchip.system.DefaultRV32Config.fir@210312.6]
  wire  _T_1792; // @[Monitor.scala 668:15:freechips.rocketchip.system.DefaultRV32Config.fir@210313.6]
  wire  _T_1794; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210315.6]
  wire  _T_1795; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210316.6]
  wire [7:0] a_size_lookup; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@210192.4 :freechips.rocketchip.system.DefaultRV32Config.fir@210193.4 Monitor.scala 633:19:freechips.rocketchip.system.DefaultRV32Config.fir@210202.4]
  wire [7:0] _GEN_86; // @[Monitor.scala 670:34:freechips.rocketchip.system.DefaultRV32Config.fir@210321.6]
  wire  _T_1796; // @[Monitor.scala 670:34:freechips.rocketchip.system.DefaultRV32Config.fir@210321.6]
  wire  _T_1798; // @[Monitor.scala 670:72:freechips.rocketchip.system.DefaultRV32Config.fir@210323.6]
  wire  _T_1799; // @[Monitor.scala 670:53:freechips.rocketchip.system.DefaultRV32Config.fir@210324.6]
  wire  _T_1801; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210326.6]
  wire  _T_1802; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210327.6]
  wire  _T_1804; // @[Monitor.scala 672:36:freechips.rocketchip.system.DefaultRV32Config.fir@210334.4]
  wire  _T_1805; // @[Monitor.scala 672:47:freechips.rocketchip.system.DefaultRV32Config.fir@210335.4]
  wire  _T_1807; // @[Monitor.scala 672:65:freechips.rocketchip.system.DefaultRV32Config.fir@210337.4]
  wire  _T_1809; // @[Monitor.scala 672:116:freechips.rocketchip.system.DefaultRV32Config.fir@210339.4]
  wire  _T_1810; // @[Monitor.scala 673:15:freechips.rocketchip.system.DefaultRV32Config.fir@210341.6]
  wire  _T_1811; // @[Monitor.scala 673:32:freechips.rocketchip.system.DefaultRV32Config.fir@210342.6]
  wire  _T_1813; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210344.6]
  wire  _T_1814; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210345.6]
  wire [2:0] a_set; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@210175.4 :freechips.rocketchip.system.DefaultRV32Config.fir@210176.4 Monitor.scala 644:13:freechips.rocketchip.system.DefaultRV32Config.fir@210230.6]
  wire [2:0] d_clr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@210254.4 :freechips.rocketchip.system.DefaultRV32Config.fir@210255.4 Monitor.scala 661:13:freechips.rocketchip.system.DefaultRV32Config.fir@210268.6]
  wire  _T_1815; // @[Monitor.scala 677:20:freechips.rocketchip.system.DefaultRV32Config.fir@210351.4]
  wire  _T_1816; // @[Monitor.scala 677:40:freechips.rocketchip.system.DefaultRV32Config.fir@210352.4]
  wire  _T_1817; // @[Monitor.scala 677:33:freechips.rocketchip.system.DefaultRV32Config.fir@210353.4]
  wire  _T_1818; // @[Monitor.scala 677:30:freechips.rocketchip.system.DefaultRV32Config.fir@210354.4]
  wire  _T_1820; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210356.4]
  wire  _T_1821; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210357.4]
  wire [2:0] _T_1822; // @[Monitor.scala 680:27:freechips.rocketchip.system.DefaultRV32Config.fir@210362.4]
  wire [2:0] _T_1823; // @[Monitor.scala 680:38:freechips.rocketchip.system.DefaultRV32Config.fir@210363.4]
  wire [2:0] _T_1824; // @[Monitor.scala 680:36:freechips.rocketchip.system.DefaultRV32Config.fir@210364.4]
  wire [11:0] a_opcodes_set; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@210177.4 :freechips.rocketchip.system.DefaultRV32Config.fir@210178.4 Monitor.scala 647:21:freechips.rocketchip.system.DefaultRV32Config.fir@210239.6]
  wire [11:0] _T_1825; // @[Monitor.scala 681:43:freechips.rocketchip.system.DefaultRV32Config.fir@210366.4]
  wire [11:0] d_opcodes_clr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@210256.4 :freechips.rocketchip.system.DefaultRV32Config.fir@210257.4 Monitor.scala 662:21:freechips.rocketchip.system.DefaultRV32Config.fir@210275.6]
  wire [11:0] _T_1826; // @[Monitor.scala 681:62:freechips.rocketchip.system.DefaultRV32Config.fir@210367.4]
  wire [11:0] _T_1827; // @[Monitor.scala 681:60:freechips.rocketchip.system.DefaultRV32Config.fir@210368.4]
  wire [23:0] a_sizes_set; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@210179.4 :freechips.rocketchip.system.DefaultRV32Config.fir@210180.4 Monitor.scala 648:19:freechips.rocketchip.system.DefaultRV32Config.fir@210242.6]
  wire [23:0] _T_1828; // @[Monitor.scala 682:39:freechips.rocketchip.system.DefaultRV32Config.fir@210370.4]
  wire [23:0] d_sizes_clr; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@210258.4 :freechips.rocketchip.system.DefaultRV32Config.fir@210259.4 Monitor.scala 663:19:freechips.rocketchip.system.DefaultRV32Config.fir@210282.6]
  wire [23:0] _T_1829; // @[Monitor.scala 682:56:freechips.rocketchip.system.DefaultRV32Config.fir@210371.4]
  wire [23:0] _T_1830; // @[Monitor.scala 682:54:freechips.rocketchip.system.DefaultRV32Config.fir@210372.4]
  reg [31:0] _T_1831; // @[Monitor.scala 684:27:freechips.rocketchip.system.DefaultRV32Config.fir@210374.4]
  wire  _T_1832; // @[Monitor.scala 687:26:freechips.rocketchip.system.DefaultRV32Config.fir@210377.4]
  wire  _T_1833; // @[Monitor.scala 687:16:freechips.rocketchip.system.DefaultRV32Config.fir@210378.4]
  wire  _T_1834; // @[Monitor.scala 687:39:freechips.rocketchip.system.DefaultRV32Config.fir@210379.4]
  wire  _T_1835; // @[Monitor.scala 687:30:freechips.rocketchip.system.DefaultRV32Config.fir@210380.4]
  wire  _T_1836; // @[Monitor.scala 687:59:freechips.rocketchip.system.DefaultRV32Config.fir@210381.4]
  wire  _T_1837; // @[Monitor.scala 687:47:freechips.rocketchip.system.DefaultRV32Config.fir@210382.4]
  wire  _T_1839; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210384.4]
  wire  _T_1840; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210385.4]
  wire [31:0] _T_1842; // @[Monitor.scala 689:26:freechips.rocketchip.system.DefaultRV32Config.fir@210391.4]
  wire  _T_1845; // @[Monitor.scala 690:27:freechips.rocketchip.system.DefaultRV32Config.fir@210395.4]
  reg [3:0] _T_1846; // @[Monitor.scala 694:27:freechips.rocketchip.system.DefaultRV32Config.fir@210399.4]
  reg [9:0] _T_1855; // @[Edges.scala 230:27:freechips.rocketchip.system.DefaultRV32Config.fir@210408.4]
  wire [9:0] _T_1857; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@210410.4]
  wire  _T_1858; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@210411.4]
  wire  _T_1868; // @[Monitor.scala 700:27:freechips.rocketchip.system.DefaultRV32Config.fir@210425.4]
  wire  _T_1871; // @[Edges.scala 72:43:freechips.rocketchip.system.DefaultRV32Config.fir@210428.4]
  wire  _T_1872; // @[Edges.scala 72:40:freechips.rocketchip.system.DefaultRV32Config.fir@210429.4]
  wire  _T_1873; // @[Monitor.scala 700:38:freechips.rocketchip.system.DefaultRV32Config.fir@210430.4]
  wire [3:0] _T_1874; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@210432.6]
  wire [3:0] _T_1875; // @[Monitor.scala 702:23:freechips.rocketchip.system.DefaultRV32Config.fir@210434.6]
  wire  _T_1877; // @[Monitor.scala 702:14:freechips.rocketchip.system.DefaultRV32Config.fir@210436.6]
  wire  _T_1879; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210438.6]
  wire  _T_1880; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210439.6]
  wire [3:0] _GEN_69; // @[Monitor.scala 700:72:freechips.rocketchip.system.DefaultRV32Config.fir@210431.4]
  wire  _T_1882; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@210447.4]
  wire [3:0] _T_1885; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@210451.6]
  wire [3:0] _T_1886; // @[Monitor.scala 708:24:freechips.rocketchip.system.DefaultRV32Config.fir@210453.6]
  wire [3:0] _T_1887; // @[Monitor.scala 708:35:freechips.rocketchip.system.DefaultRV32Config.fir@210454.6]
  wire  _T_1890; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210457.6]
  wire  _T_1891; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210458.6]
  wire [3:0] _GEN_70; // @[Monitor.scala 706:73:freechips.rocketchip.system.DefaultRV32Config.fir@210450.4]
  wire [3:0] _T_1892; // @[Monitor.scala 713:27:freechips.rocketchip.system.DefaultRV32Config.fir@210464.4]
  wire [3:0] _T_1893; // @[Monitor.scala 713:38:freechips.rocketchip.system.DefaultRV32Config.fir@210465.4]
  wire [3:0] _T_1894; // @[Monitor.scala 713:36:freechips.rocketchip.system.DefaultRV32Config.fir@210466.4]
  wire  _GEN_87; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207660.10]
  wire  _GEN_103; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207789.10]
  wire  _GEN_121; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207929.10]
  wire  _GEN_133; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208036.10]
  wire  _GEN_143; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208135.10]
  wire  _GEN_153; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208226.10]
  wire  _GEN_163; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208315.10]
  wire  _GEN_173; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208404.10]
  wire  _GEN_185; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208473.10]
  wire  _GEN_195; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208515.10]
  wire  _GEN_205; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208573.10]
  wire  _GEN_215; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208632.10]
  wire  _GEN_221; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208667.10]
  wire  _GEN_227; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208703.10]
  wire  _GEN_233; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208902.10]
  wire  _GEN_247; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208957.10]
  wire  _GEN_261; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209012.10]
  wire  _GEN_273; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209059.10]
  wire  _GEN_285; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209108.10]
  wire  _GEN_295; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209155.10]
  wire  _GEN_305; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209202.10]
  wire  _GEN_317; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209358.10]
  wire  _GEN_327; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209406.10]
  wire  _GEN_337; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209495.10]
  wire  _GEN_349; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209615.10]
  wire  _GEN_361; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209678.10]
  wire  _GEN_369; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209718.10]
  wire  _GEN_377; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209750.10]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11:freechips.rocketchip.system.DefaultRV32Config.fir@210375.4]
    .out(plusarg_reader_out)
  );
  assign _T_4 = io_in_a_bits_source == 2'h0; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@207523.6]
  assign _T_5 = io_in_a_bits_source == 2'h1; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@207524.6]
  assign _T_6 = io_in_a_bits_source == 2'h2; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@207525.6]
  assign _T_8 = _T_4 | _T_5; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@207531.6]
  assign _T_9 = _T_8 | _T_6; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@207532.6]
  assign _T_11 = 27'hfff << io_in_a_bits_size; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@207534.6]
  assign _T_13 = ~_T_11[11:0]; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@207536.6]
  assign _GEN_71 = {{20'd0}, _T_13}; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@207537.6]
  assign _T_14 = io_in_a_bits_address & _GEN_71; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@207537.6]
  assign _T_15 = _T_14 == 32'h0; // @[Edges.scala 22:24:freechips.rocketchip.system.DefaultRV32Config.fir@207538.6]
  assign _T_18 = 2'h1 << io_in_a_bits_size[0]; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@207541.6]
  assign _T_20 = _T_18 | 2'h1; // @[Misc.scala 201:81:freechips.rocketchip.system.DefaultRV32Config.fir@207543.6]
  assign _T_21 = io_in_a_bits_size >= 4'h2; // @[Misc.scala 205:21:freechips.rocketchip.system.DefaultRV32Config.fir@207544.6]
  assign _T_24 = ~io_in_a_bits_address[1]; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@207547.6]
  assign _T_26 = _T_20[1] & _T_24; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@207549.6]
  assign _T_27 = _T_21 | _T_26; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@207550.6]
  assign _T_29 = _T_20[1] & io_in_a_bits_address[1]; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@207552.6]
  assign _T_30 = _T_21 | _T_29; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@207553.6]
  assign _T_33 = ~io_in_a_bits_address[0]; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@207556.6]
  assign _T_34 = _T_24 & _T_33; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@207557.6]
  assign _T_35 = _T_20[0] & _T_34; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@207558.6]
  assign _T_36 = _T_27 | _T_35; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@207559.6]
  assign _T_37 = _T_24 & io_in_a_bits_address[0]; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@207560.6]
  assign _T_38 = _T_20[0] & _T_37; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@207561.6]
  assign _T_39 = _T_27 | _T_38; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@207562.6]
  assign _T_40 = io_in_a_bits_address[1] & _T_33; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@207563.6]
  assign _T_41 = _T_20[0] & _T_40; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@207564.6]
  assign _T_42 = _T_30 | _T_41; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@207565.6]
  assign _T_43 = io_in_a_bits_address[1] & io_in_a_bits_address[0]; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@207566.6]
  assign _T_44 = _T_20[0] & _T_43; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@207567.6]
  assign _T_45 = _T_30 | _T_44; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@207568.6]
  assign _T_48 = {_T_45,_T_42,_T_39,_T_36}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@207571.6]
  assign _T_52 = {1'b0,$signed(io_in_a_bits_address)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@207575.6]
  assign _T_78 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 79:25:freechips.rocketchip.system.DefaultRV32Config.fir@207605.6]
  assign _T_83 = $signed(_T_52) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@207611.8]
  assign _T_84 = $signed(_T_83) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@207612.8]
  assign _T_85 = io_in_a_bits_address ^ 32'h3000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@207613.8]
  assign _T_86 = {1'b0,$signed(_T_85)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@207614.8]
  assign _T_88 = $signed(_T_86) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@207616.8]
  assign _T_89 = $signed(_T_88) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@207617.8]
  assign _T_90 = io_in_a_bits_address ^ 32'h10000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@207618.8]
  assign _T_91 = {1'b0,$signed(_T_90)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@207619.8]
  assign _T_93 = $signed(_T_91) & -33'sh10000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@207621.8]
  assign _T_94 = $signed(_T_93) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@207622.8]
  assign _T_95 = io_in_a_bits_address ^ 32'h2000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@207623.8]
  assign _T_96 = {1'b0,$signed(_T_95)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@207624.8]
  assign _T_98 = $signed(_T_96) & -33'sh10000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@207626.8]
  assign _T_99 = $signed(_T_98) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@207627.8]
  assign _T_100 = io_in_a_bits_address ^ 32'hc000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@207628.8]
  assign _T_101 = {1'b0,$signed(_T_100)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@207629.8]
  assign _T_103 = $signed(_T_101) & -33'sh4000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@207631.8]
  assign _T_104 = $signed(_T_103) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@207632.8]
  assign _T_105 = io_in_a_bits_address ^ 32'h60000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@207633.8]
  assign _T_106 = {1'b0,$signed(_T_105)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@207634.8]
  assign _T_108 = $signed(_T_106) & -33'sh20000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@207636.8]
  assign _T_109 = $signed(_T_108) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@207637.8]
  assign _T_110 = _T_84 | _T_89; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@207638.8]
  assign _T_117 = io_in_a_bits_size <= 4'h6; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@207645.8]
  assign _T_120 = io_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@207648.8]
  assign _T_121 = {1'b0,$signed(_T_120)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@207649.8]
  assign _T_123 = $signed(_T_121) & -33'sh10000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@207651.8]
  assign _T_124 = $signed(_T_123) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@207652.8]
  assign _T_125 = _T_117 & _T_124; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@207653.8]
  assign _T_129 = _T_125 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207657.8]
  assign _T_130 = ~_T_129; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207658.8]
  assign _T_135 = 4'h6 == io_in_a_bits_size; // @[Parameters.scala 92:48:freechips.rocketchip.system.DefaultRV32Config.fir@207671.8]
  assign _T_136 = _T_4 & _T_135; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@207672.8]
  assign _T_143 = _T_136 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207680.8]
  assign _T_144 = ~_T_143; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207681.8]
  assign _T_146 = _T_9 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207687.8]
  assign _T_147 = ~_T_146; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207688.8]
  assign _T_150 = _T_21 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207695.8]
  assign _T_151 = ~_T_150; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207696.8]
  assign _T_153 = _T_15 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207702.8]
  assign _T_154 = ~_T_153; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207703.8]
  assign _T_155 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 110:27:freechips.rocketchip.system.DefaultRV32Config.fir@207708.8]
  assign _T_157 = _T_155 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207710.8]
  assign _T_158 = ~_T_157; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207711.8]
  assign _T_159 = ~io_in_a_bits_mask; // @[Monitor.scala 86:18:freechips.rocketchip.system.DefaultRV32Config.fir@207716.8]
  assign _T_160 = _T_159 == 4'h0; // @[Monitor.scala 86:31:freechips.rocketchip.system.DefaultRV32Config.fir@207717.8]
  assign _T_162 = _T_160 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207719.8]
  assign _T_163 = ~_T_162; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207720.8]
  assign _T_164 = ~io_in_a_bits_corrupt; // @[Monitor.scala 87:18:freechips.rocketchip.system.DefaultRV32Config.fir@207725.8]
  assign _T_166 = _T_164 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207727.8]
  assign _T_167 = ~_T_166; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207728.8]
  assign _T_168 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 90:25:freechips.rocketchip.system.DefaultRV32Config.fir@207734.6]
  assign _T_249 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 97:31:freechips.rocketchip.system.DefaultRV32Config.fir@207845.8]
  assign _T_251 = _T_249 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207847.8]
  assign _T_252 = ~_T_251; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207848.8]
  assign _T_262 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 102:25:freechips.rocketchip.system.DefaultRV32Config.fir@207871.6]
  assign _T_264 = io_in_a_bits_size <= 4'hc; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@207874.8]
  assign _T_272 = _T_264 & _T_89; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@207882.8]
  assign _T_307 = _T_84 | _T_94; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@207917.8]
  assign _T_308 = _T_307 | _T_99; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@207918.8]
  assign _T_309 = _T_308 | _T_104; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@207919.8]
  assign _T_310 = _T_309 | _T_109; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@207920.8]
  assign _T_311 = _T_310 | _T_124; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@207921.8]
  assign _T_312 = _T_117 & _T_311; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@207922.8]
  assign _T_314 = _T_272 | _T_312; // @[Parameters.scala 553:30:freechips.rocketchip.system.DefaultRV32Config.fir@207924.8]
  assign _T_316 = _T_314 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207926.8]
  assign _T_317 = ~_T_316; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207927.8]
  assign _T_324 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 106:31:freechips.rocketchip.system.DefaultRV32Config.fir@207946.8]
  assign _T_326 = _T_324 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207948.8]
  assign _T_327 = ~_T_326; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207949.8]
  assign _T_328 = io_in_a_bits_mask == _T_48; // @[Monitor.scala 107:30:freechips.rocketchip.system.DefaultRV32Config.fir@207954.8]
  assign _T_330 = _T_328 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207956.8]
  assign _T_331 = ~_T_330; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207957.8]
  assign _T_336 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 111:25:freechips.rocketchip.system.DefaultRV32Config.fir@207971.6]
  assign _T_371 = _T_84 | _T_99; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@208007.8]
  assign _T_372 = _T_371 | _T_104; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@208008.8]
  assign _T_373 = _T_372 | _T_124; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@208009.8]
  assign _T_374 = _T_117 & _T_373; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@208010.8]
  assign _T_383 = io_in_a_bits_size <= 4'h8; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@208019.8]
  assign _T_391 = _T_383 & _T_109; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@208027.8]
  assign _T_393 = _T_272 | _T_374; // @[Parameters.scala 553:30:freechips.rocketchip.system.DefaultRV32Config.fir@208029.8]
  assign _T_395 = _T_393 | _T_391; // @[Parameters.scala 553:30:freechips.rocketchip.system.DefaultRV32Config.fir@208031.8]
  assign _T_397 = _T_395 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208033.8]
  assign _T_398 = ~_T_397; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208034.8]
  assign _T_413 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 119:25:freechips.rocketchip.system.DefaultRV32Config.fir@208070.6]
  assign _T_486 = ~_T_48; // @[Monitor.scala 124:33:freechips.rocketchip.system.DefaultRV32Config.fir@208160.8]
  assign _T_487 = io_in_a_bits_mask & _T_486; // @[Monitor.scala 124:31:freechips.rocketchip.system.DefaultRV32Config.fir@208161.8]
  assign _T_488 = _T_487 == 4'h0; // @[Monitor.scala 124:40:freechips.rocketchip.system.DefaultRV32Config.fir@208162.8]
  assign _T_490 = _T_488 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208164.8]
  assign _T_491 = ~_T_490; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208165.8]
  assign _T_492 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 127:25:freechips.rocketchip.system.DefaultRV32Config.fir@208171.6]
  assign _T_494 = io_in_a_bits_size <= 4'h2; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@208174.8]
  assign _T_518 = _T_110 | _T_99; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@208198.8]
  assign _T_519 = _T_518 | _T_104; // @[Parameters.scala 552:42:freechips.rocketchip.system.DefaultRV32Config.fir@208199.8]
  assign _T_520 = _T_494 & _T_519; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@208200.8]
  assign _T_543 = _T_520 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208223.8]
  assign _T_544 = ~_T_543; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208224.8]
  assign _T_551 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 140:33:freechips.rocketchip.system.DefaultRV32Config.fir@208243.8]
  assign _T_553 = _T_551 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208245.8]
  assign _T_554 = ~_T_553; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208246.8]
  assign _T_559 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 135:25:freechips.rocketchip.system.DefaultRV32Config.fir@208260.6]
  assign _T_618 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 147:30:freechips.rocketchip.system.DefaultRV32Config.fir@208332.8]
  assign _T_620 = _T_618 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208334.8]
  assign _T_621 = ~_T_620; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208335.8]
  assign _T_626 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 143:25:freechips.rocketchip.system.DefaultRV32Config.fir@208349.6]
  assign _T_677 = _T_272 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208401.8]
  assign _T_678 = ~_T_677; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208402.8]
  assign _T_685 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 160:28:freechips.rocketchip.system.DefaultRV32Config.fir@208421.8]
  assign _T_687 = _T_685 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208423.8]
  assign _T_688 = ~_T_687; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208424.8]
  assign _T_697 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 44:24:freechips.rocketchip.system.DefaultRV32Config.fir@208448.6]
  assign _T_699 = _T_697 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208450.6]
  assign _T_700 = ~_T_699; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208451.6]
  assign _T_701 = io_in_d_bits_source == 2'h0; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@208456.6]
  assign _T_702 = io_in_d_bits_source == 2'h1; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@208457.6]
  assign _T_703 = io_in_d_bits_source == 2'h2; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@208458.6]
  assign _T_705 = _T_701 | _T_702; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@208464.6]
  assign _T_706 = _T_705 | _T_703; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@208465.6]
  assign _T_708 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 307:25:freechips.rocketchip.system.DefaultRV32Config.fir@208467.6]
  assign _T_710 = _T_706 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208470.8]
  assign _T_711 = ~_T_710; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208471.8]
  assign _T_712 = io_in_d_bits_size >= 4'h2; // @[Monitor.scala 309:27:freechips.rocketchip.system.DefaultRV32Config.fir@208476.8]
  assign _T_714 = _T_712 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208478.8]
  assign _T_715 = ~_T_714; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208479.8]
  assign _T_716 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 310:28:freechips.rocketchip.system.DefaultRV32Config.fir@208484.8]
  assign _T_718 = _T_716 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208486.8]
  assign _T_719 = ~_T_718; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208487.8]
  assign _T_720 = ~io_in_d_bits_corrupt; // @[Monitor.scala 311:15:freechips.rocketchip.system.DefaultRV32Config.fir@208492.8]
  assign _T_722 = _T_720 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208494.8]
  assign _T_723 = ~_T_722; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208495.8]
  assign _T_724 = ~io_in_d_bits_denied; // @[Monitor.scala 312:15:freechips.rocketchip.system.DefaultRV32Config.fir@208500.8]
  assign _T_726 = _T_724 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208502.8]
  assign _T_727 = ~_T_726; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208503.8]
  assign _T_728 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 315:25:freechips.rocketchip.system.DefaultRV32Config.fir@208509.6]
  assign _T_739 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 104:26:freechips.rocketchip.system.DefaultRV32Config.fir@208533.8]
  assign _T_741 = _T_739 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208535.8]
  assign _T_742 = ~_T_741; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208536.8]
  assign _T_743 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 320:28:freechips.rocketchip.system.DefaultRV32Config.fir@208541.8]
  assign _T_745 = _T_743 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208543.8]
  assign _T_746 = ~_T_745; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208544.8]
  assign _T_756 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 325:25:freechips.rocketchip.system.DefaultRV32Config.fir@208567.6]
  assign _T_776 = _T_724 | io_in_d_bits_corrupt; // @[Monitor.scala 331:30:freechips.rocketchip.system.DefaultRV32Config.fir@208608.8]
  assign _T_778 = _T_776 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208610.8]
  assign _T_779 = ~_T_778; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208611.8]
  assign _T_785 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 335:25:freechips.rocketchip.system.DefaultRV32Config.fir@208626.6]
  assign _T_802 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 343:25:freechips.rocketchip.system.DefaultRV32Config.fir@208661.6]
  assign _T_820 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 351:25:freechips.rocketchip.system.DefaultRV32Config.fir@208697.6]
  assign _T_837 = io_in_b_bits_opcode <= 3'h6; // @[Bundles.scala 42:24:freechips.rocketchip.system.DefaultRV32Config.fir@208734.6]
  assign _T_839 = _T_837 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208736.6]
  assign _T_840 = ~_T_839; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208737.6]
  assign _T_841 = io_in_b_bits_source == 2'h0; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@208742.6]
  assign _T_844 = {1'b0,$signed(io_in_b_bits_address)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208745.6]
  assign _T_849 = io_in_b_bits_source == 2'h1; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@208750.6]
  assign _T_857 = io_in_b_bits_source == 2'h2; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@208758.6]
  assign _T_870 = io_in_b_bits_address ^ 32'h3000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@208775.6]
  assign _T_871 = {1'b0,$signed(_T_870)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208776.6]
  assign _T_873 = $signed(_T_871) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208778.6]
  assign _T_874 = $signed(_T_873) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208779.6]
  assign _T_875 = io_in_b_bits_address ^ 32'hc000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@208780.6]
  assign _T_876 = {1'b0,$signed(_T_875)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208781.6]
  assign _T_878 = $signed(_T_876) & -33'sh4000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208783.6]
  assign _T_879 = $signed(_T_878) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208784.6]
  assign _T_880 = io_in_b_bits_address ^ 32'h2000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@208785.6]
  assign _T_881 = {1'b0,$signed(_T_880)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208786.6]
  assign _T_883 = $signed(_T_881) & -33'sh10000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208788.6]
  assign _T_884 = $signed(_T_883) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208789.6]
  assign _T_888 = $signed(_T_844) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208793.6]
  assign _T_889 = $signed(_T_888) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208794.6]
  assign _T_890 = io_in_b_bits_address ^ 32'h10000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@208795.6]
  assign _T_891 = {1'b0,$signed(_T_890)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208796.6]
  assign _T_893 = $signed(_T_891) & -33'sh10000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208798.6]
  assign _T_894 = $signed(_T_893) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208799.6]
  assign _T_895 = io_in_b_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@208800.6]
  assign _T_896 = {1'b0,$signed(_T_895)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208801.6]
  assign _T_898 = $signed(_T_896) & -33'sh10000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208803.6]
  assign _T_899 = $signed(_T_898) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208804.6]
  assign _T_900 = io_in_b_bits_address ^ 32'h60000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@208805.6]
  assign _T_901 = {1'b0,$signed(_T_900)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@208806.6]
  assign _T_903 = $signed(_T_901) & -33'sh20000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@208808.6]
  assign _T_904 = $signed(_T_903) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@208809.6]
  assign _T_906 = _T_874 | _T_879; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@208819.6]
  assign _T_907 = _T_906 | _T_884; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@208820.6]
  assign _T_908 = _T_907 | _T_889; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@208821.6]
  assign _T_909 = _T_908 | _T_894; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@208822.6]
  assign _T_910 = _T_909 | _T_899; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@208823.6]
  assign _T_911 = _T_910 | _T_904; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@208824.6]
  assign _T_913 = 27'hfff << io_in_b_bits_size; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@208826.6]
  assign _T_915 = ~_T_913[11:0]; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@208828.6]
  assign _GEN_72 = {{20'd0}, _T_915}; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@208829.6]
  assign _T_916 = io_in_b_bits_address & _GEN_72; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@208829.6]
  assign _T_917 = _T_916 == 32'h0; // @[Edges.scala 22:24:freechips.rocketchip.system.DefaultRV32Config.fir@208830.6]
  assign _T_920 = 2'h1 << io_in_b_bits_size[0]; // @[OneHot.scala 65:12:freechips.rocketchip.system.DefaultRV32Config.fir@208833.6]
  assign _T_922 = _T_920 | 2'h1; // @[Misc.scala 201:81:freechips.rocketchip.system.DefaultRV32Config.fir@208835.6]
  assign _T_923 = io_in_b_bits_size >= 4'h2; // @[Misc.scala 205:21:freechips.rocketchip.system.DefaultRV32Config.fir@208836.6]
  assign _T_926 = ~io_in_b_bits_address[1]; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@208839.6]
  assign _T_928 = _T_922[1] & _T_926; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@208841.6]
  assign _T_929 = _T_923 | _T_928; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@208842.6]
  assign _T_931 = _T_922[1] & io_in_b_bits_address[1]; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@208844.6]
  assign _T_932 = _T_923 | _T_931; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@208845.6]
  assign _T_935 = ~io_in_b_bits_address[0]; // @[Misc.scala 210:20:freechips.rocketchip.system.DefaultRV32Config.fir@208848.6]
  assign _T_936 = _T_926 & _T_935; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@208849.6]
  assign _T_937 = _T_922[0] & _T_936; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@208850.6]
  assign _T_938 = _T_929 | _T_937; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@208851.6]
  assign _T_939 = _T_926 & io_in_b_bits_address[0]; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@208852.6]
  assign _T_940 = _T_922[0] & _T_939; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@208853.6]
  assign _T_941 = _T_929 | _T_940; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@208854.6]
  assign _T_942 = io_in_b_bits_address[1] & _T_935; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@208855.6]
  assign _T_943 = _T_922[0] & _T_942; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@208856.6]
  assign _T_944 = _T_932 | _T_943; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@208857.6]
  assign _T_945 = io_in_b_bits_address[1] & io_in_b_bits_address[0]; // @[Misc.scala 213:27:freechips.rocketchip.system.DefaultRV32Config.fir@208858.6]
  assign _T_946 = _T_922[0] & _T_945; // @[Misc.scala 214:38:freechips.rocketchip.system.DefaultRV32Config.fir@208859.6]
  assign _T_947 = _T_932 | _T_946; // @[Misc.scala 214:29:freechips.rocketchip.system.DefaultRV32Config.fir@208860.6]
  assign _T_950 = {_T_947,_T_944,_T_941,_T_938}; // @[Cat.scala 29:58:freechips.rocketchip.system.DefaultRV32Config.fir@208863.6]
  assign _T_957 = _T_857 ? 2'h2 : 2'h0; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@208874.6]
  assign _GEN_73 = {{1'd0}, _T_849}; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@208876.6]
  assign _T_959 = _GEN_73 | _T_957; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@208876.6]
  assign _T_961 = _T_959 == io_in_b_bits_source; // @[Monitor.scala 162:113:freechips.rocketchip.system.DefaultRV32Config.fir@208879.6]
  assign _T_962 = io_in_b_bits_opcode == 3'h6; // @[Monitor.scala 164:25:freechips.rocketchip.system.DefaultRV32Config.fir@208880.6]
  assign _T_967 = 4'h6 == io_in_b_bits_size; // @[Parameters.scala 92:48:freechips.rocketchip.system.DefaultRV32Config.fir@208890.8]
  assign _T_968 = _T_841 & _T_967; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@208891.8]
  assign _T_975 = _T_968 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208899.8]
  assign _T_976 = ~_T_975; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208900.8]
  assign _T_978 = _T_911 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208906.8]
  assign _T_979 = ~_T_978; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208907.8]
  assign _T_981 = _T_961 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208913.8]
  assign _T_982 = ~_T_981; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208914.8]
  assign _T_984 = _T_917 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208920.8]
  assign _T_985 = ~_T_984; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208921.8]
  assign _T_986 = io_in_b_bits_param <= 2'h2; // @[Bundles.scala 104:26:freechips.rocketchip.system.DefaultRV32Config.fir@208926.8]
  assign _T_988 = _T_986 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208928.8]
  assign _T_989 = ~_T_988; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208929.8]
  assign _T_990 = io_in_b_bits_mask == _T_950; // @[Monitor.scala 170:30:freechips.rocketchip.system.DefaultRV32Config.fir@208934.8]
  assign _T_992 = _T_990 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208936.8]
  assign _T_993 = ~_T_992; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208937.8]
  assign _T_994 = ~io_in_b_bits_corrupt; // @[Monitor.scala 171:18:freechips.rocketchip.system.DefaultRV32Config.fir@208942.8]
  assign _T_996 = _T_994 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208944.8]
  assign _T_997 = ~_T_996; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208945.8]
  assign _T_998 = io_in_b_bits_opcode == 3'h4; // @[Monitor.scala 174:25:freechips.rocketchip.system.DefaultRV32Config.fir@208951.6]
  assign _T_1001 = ~reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208955.8]
  assign _T_1011 = io_in_b_bits_param == 2'h0; // @[Monitor.scala 179:31:freechips.rocketchip.system.DefaultRV32Config.fir@208981.8]
  assign _T_1013 = _T_1011 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208983.8]
  assign _T_1014 = ~_T_1013; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208984.8]
  assign _T_1023 = io_in_b_bits_opcode == 3'h0; // @[Monitor.scala 184:25:freechips.rocketchip.system.DefaultRV32Config.fir@209006.6]
  assign _T_1044 = io_in_b_bits_opcode == 3'h1; // @[Monitor.scala 193:25:freechips.rocketchip.system.DefaultRV32Config.fir@209053.6]
  assign _T_1061 = ~_T_950; // @[Monitor.scala 199:33:freechips.rocketchip.system.DefaultRV32Config.fir@209091.8]
  assign _T_1062 = io_in_b_bits_mask & _T_1061; // @[Monitor.scala 199:31:freechips.rocketchip.system.DefaultRV32Config.fir@209092.8]
  assign _T_1063 = _T_1062 == 4'h0; // @[Monitor.scala 199:40:freechips.rocketchip.system.DefaultRV32Config.fir@209093.8]
  assign _T_1065 = _T_1063 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209095.8]
  assign _T_1066 = ~_T_1065; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209096.8]
  assign _T_1067 = io_in_b_bits_opcode == 3'h2; // @[Monitor.scala 202:25:freechips.rocketchip.system.DefaultRV32Config.fir@209102.6]
  assign _T_1088 = io_in_b_bits_opcode == 3'h3; // @[Monitor.scala 211:25:freechips.rocketchip.system.DefaultRV32Config.fir@209149.6]
  assign _T_1109 = io_in_b_bits_opcode == 3'h5; // @[Monitor.scala 220:25:freechips.rocketchip.system.DefaultRV32Config.fir@209196.6]
  assign _T_1134 = io_in_c_bits_source == 2'h0; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@209253.6]
  assign _T_1135 = io_in_c_bits_source == 2'h1; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@209254.6]
  assign _T_1136 = io_in_c_bits_source == 2'h2; // @[Parameters.scala 47:9:freechips.rocketchip.system.DefaultRV32Config.fir@209255.6]
  assign _T_1138 = _T_1134 | _T_1135; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@209261.6]
  assign _T_1139 = _T_1138 | _T_1136; // @[Parameters.scala 924:46:freechips.rocketchip.system.DefaultRV32Config.fir@209262.6]
  assign _T_1141 = 27'hfff << io_in_c_bits_size; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@209264.6]
  assign _T_1143 = ~_T_1141[11:0]; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@209266.6]
  assign _GEN_74 = {{20'd0}, _T_1143}; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@209267.6]
  assign _T_1144 = io_in_c_bits_address & _GEN_74; // @[Edges.scala 22:16:freechips.rocketchip.system.DefaultRV32Config.fir@209267.6]
  assign _T_1145 = _T_1144 == 32'h0; // @[Edges.scala 22:24:freechips.rocketchip.system.DefaultRV32Config.fir@209268.6]
  assign _T_1146 = io_in_c_bits_address ^ 32'h3000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@209269.6]
  assign _T_1147 = {1'b0,$signed(_T_1146)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@209270.6]
  assign _T_1149 = $signed(_T_1147) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@209272.6]
  assign _T_1150 = $signed(_T_1149) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@209273.6]
  assign _T_1151 = io_in_c_bits_address ^ 32'hc000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@209274.6]
  assign _T_1152 = {1'b0,$signed(_T_1151)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@209275.6]
  assign _T_1154 = $signed(_T_1152) & -33'sh4000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@209277.6]
  assign _T_1155 = $signed(_T_1154) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@209278.6]
  assign _T_1156 = io_in_c_bits_address ^ 32'h2000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@209279.6]
  assign _T_1157 = {1'b0,$signed(_T_1156)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@209280.6]
  assign _T_1159 = $signed(_T_1157) & -33'sh10000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@209282.6]
  assign _T_1160 = $signed(_T_1159) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@209283.6]
  assign _T_1162 = {1'b0,$signed(io_in_c_bits_address)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@209285.6]
  assign _T_1164 = $signed(_T_1162) & -33'sh1000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@209287.6]
  assign _T_1165 = $signed(_T_1164) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@209288.6]
  assign _T_1166 = io_in_c_bits_address ^ 32'h10000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@209289.6]
  assign _T_1167 = {1'b0,$signed(_T_1166)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@209290.6]
  assign _T_1169 = $signed(_T_1167) & -33'sh10000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@209292.6]
  assign _T_1170 = $signed(_T_1169) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@209293.6]
  assign _T_1171 = io_in_c_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@209294.6]
  assign _T_1172 = {1'b0,$signed(_T_1171)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@209295.6]
  assign _T_1174 = $signed(_T_1172) & -33'sh10000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@209297.6]
  assign _T_1175 = $signed(_T_1174) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@209298.6]
  assign _T_1176 = io_in_c_bits_address ^ 32'h60000000; // @[Parameters.scala 137:31:freechips.rocketchip.system.DefaultRV32Config.fir@209299.6]
  assign _T_1177 = {1'b0,$signed(_T_1176)}; // @[Parameters.scala 137:49:freechips.rocketchip.system.DefaultRV32Config.fir@209300.6]
  assign _T_1179 = $signed(_T_1177) & -33'sh20000000; // @[Parameters.scala 137:52:freechips.rocketchip.system.DefaultRV32Config.fir@209302.6]
  assign _T_1180 = $signed(_T_1179) == 33'sh0; // @[Parameters.scala 137:67:freechips.rocketchip.system.DefaultRV32Config.fir@209303.6]
  assign _T_1182 = _T_1150 | _T_1155; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@209313.6]
  assign _T_1183 = _T_1182 | _T_1160; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@209314.6]
  assign _T_1184 = _T_1183 | _T_1165; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@209315.6]
  assign _T_1185 = _T_1184 | _T_1170; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@209316.6]
  assign _T_1186 = _T_1185 | _T_1175; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@209317.6]
  assign _T_1187 = _T_1186 | _T_1180; // @[Parameters.scala 535:64:freechips.rocketchip.system.DefaultRV32Config.fir@209318.6]
  assign _T_1217 = io_in_c_bits_opcode == 3'h4; // @[Monitor.scala 239:25:freechips.rocketchip.system.DefaultRV32Config.fir@209352.6]
  assign _T_1219 = _T_1187 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209355.8]
  assign _T_1220 = ~_T_1219; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209356.8]
  assign _T_1222 = _T_1139 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209362.8]
  assign _T_1223 = ~_T_1222; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209363.8]
  assign _T_1224 = io_in_c_bits_size >= 4'h2; // @[Monitor.scala 242:30:freechips.rocketchip.system.DefaultRV32Config.fir@209368.8]
  assign _T_1226 = _T_1224 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209370.8]
  assign _T_1227 = ~_T_1226; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209371.8]
  assign _T_1229 = _T_1145 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209377.8]
  assign _T_1230 = ~_T_1229; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209378.8]
  assign _T_1231 = io_in_c_bits_param <= 3'h5; // @[Bundles.scala 122:29:freechips.rocketchip.system.DefaultRV32Config.fir@209383.8]
  assign _T_1233 = _T_1231 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209385.8]
  assign _T_1234 = ~_T_1233; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209386.8]
  assign _T_1239 = io_in_c_bits_opcode == 3'h5; // @[Monitor.scala 248:25:freechips.rocketchip.system.DefaultRV32Config.fir@209400.6]
  assign _T_1257 = io_in_c_bits_opcode == 3'h6; // @[Monitor.scala 256:25:freechips.rocketchip.system.DefaultRV32Config.fir@209440.6]
  assign _T_1296 = io_in_c_bits_size <= 4'h6; // @[Parameters.scala 93:42:freechips.rocketchip.system.DefaultRV32Config.fir@209480.8]
  assign _T_1304 = _T_1296 & _T_1175; // @[Parameters.scala 551:56:freechips.rocketchip.system.DefaultRV32Config.fir@209488.8]
  assign _T_1308 = _T_1304 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209492.8]
  assign _T_1309 = ~_T_1308; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209493.8]
  assign _T_1314 = 4'h6 == io_in_c_bits_size; // @[Parameters.scala 92:48:freechips.rocketchip.system.DefaultRV32Config.fir@209506.8]
  assign _T_1315 = _T_1134 & _T_1314; // @[Mux.scala 27:72:freechips.rocketchip.system.DefaultRV32Config.fir@209507.8]
  assign _T_1322 = _T_1315 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209515.8]
  assign _T_1323 = ~_T_1322; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209516.8]
  assign _T_1334 = io_in_c_bits_param <= 3'h2; // @[Bundles.scala 116:29:freechips.rocketchip.system.DefaultRV32Config.fir@209543.8]
  assign _T_1336 = _T_1334 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209545.8]
  assign _T_1337 = ~_T_1336; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209546.8]
  assign _T_1342 = io_in_c_bits_opcode == 3'h7; // @[Monitor.scala 266:25:freechips.rocketchip.system.DefaultRV32Config.fir@209560.6]
  assign _T_1423 = io_in_c_bits_opcode == 3'h0; // @[Monitor.scala 275:25:freechips.rocketchip.system.DefaultRV32Config.fir@209672.6]
  assign _T_1433 = io_in_c_bits_param == 3'h0; // @[Monitor.scala 279:31:freechips.rocketchip.system.DefaultRV32Config.fir@209695.8]
  assign _T_1435 = _T_1433 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209697.8]
  assign _T_1436 = ~_T_1435; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209698.8]
  assign _T_1441 = io_in_c_bits_opcode == 3'h1; // @[Monitor.scala 283:25:freechips.rocketchip.system.DefaultRV32Config.fir@209712.6]
  assign _T_1455 = io_in_c_bits_opcode == 3'h2; // @[Monitor.scala 290:25:freechips.rocketchip.system.DefaultRV32Config.fir@209744.6]
  assign _T_1477 = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@209795.4]
  assign _T_1484 = ~io_in_a_bits_opcode[2]; // @[Edges.scala 93:28:freechips.rocketchip.system.DefaultRV32Config.fir@209802.4]
  assign _T_1488 = _T_1486 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@209806.4]
  assign _T_1489 = _T_1486 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@209807.4]
  assign _T_1502 = ~_T_1489; // @[Monitor.scala 386:22:freechips.rocketchip.system.DefaultRV32Config.fir@209823.4]
  assign _T_1503 = io_in_a_valid & _T_1502; // @[Monitor.scala 386:19:freechips.rocketchip.system.DefaultRV32Config.fir@209824.4]
  assign _T_1504 = io_in_a_bits_opcode == _T_1497; // @[Monitor.scala 387:32:freechips.rocketchip.system.DefaultRV32Config.fir@209826.6]
  assign _T_1506 = _T_1504 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209828.6]
  assign _T_1507 = ~_T_1506; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209829.6]
  assign _T_1508 = io_in_a_bits_param == _T_1498; // @[Monitor.scala 388:32:freechips.rocketchip.system.DefaultRV32Config.fir@209834.6]
  assign _T_1510 = _T_1508 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209836.6]
  assign _T_1511 = ~_T_1510; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209837.6]
  assign _T_1512 = io_in_a_bits_size == _T_1499; // @[Monitor.scala 389:32:freechips.rocketchip.system.DefaultRV32Config.fir@209842.6]
  assign _T_1514 = _T_1512 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209844.6]
  assign _T_1515 = ~_T_1514; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209845.6]
  assign _T_1516 = io_in_a_bits_source == _T_1500; // @[Monitor.scala 390:32:freechips.rocketchip.system.DefaultRV32Config.fir@209850.6]
  assign _T_1518 = _T_1516 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209852.6]
  assign _T_1519 = ~_T_1518; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209853.6]
  assign _T_1520 = io_in_a_bits_address == _T_1501; // @[Monitor.scala 391:32:freechips.rocketchip.system.DefaultRV32Config.fir@209858.6]
  assign _T_1522 = _T_1520 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209860.6]
  assign _T_1523 = ~_T_1522; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209861.6]
  assign _T_1525 = _T_1477 & _T_1489; // @[Monitor.scala 393:20:freechips.rocketchip.system.DefaultRV32Config.fir@209868.4]
  assign _T_1526 = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@209876.4]
  assign _T_1528 = 27'hfff << io_in_d_bits_size; // @[package.scala 207:77:freechips.rocketchip.system.DefaultRV32Config.fir@209878.4]
  assign _T_1530 = ~_T_1528[11:0]; // @[package.scala 207:46:freechips.rocketchip.system.DefaultRV32Config.fir@209880.4]
  assign _T_1536 = _T_1534 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@209886.4]
  assign _T_1537 = _T_1534 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@209887.4]
  assign _T_1551 = ~_T_1537; // @[Monitor.scala 538:22:freechips.rocketchip.system.DefaultRV32Config.fir@209904.4]
  assign _T_1552 = io_in_d_valid & _T_1551; // @[Monitor.scala 538:19:freechips.rocketchip.system.DefaultRV32Config.fir@209905.4]
  assign _T_1553 = io_in_d_bits_opcode == _T_1545; // @[Monitor.scala 539:29:freechips.rocketchip.system.DefaultRV32Config.fir@209907.6]
  assign _T_1555 = _T_1553 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209909.6]
  assign _T_1556 = ~_T_1555; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209910.6]
  assign _T_1557 = io_in_d_bits_param == _T_1546; // @[Monitor.scala 540:29:freechips.rocketchip.system.DefaultRV32Config.fir@209915.6]
  assign _T_1559 = _T_1557 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209917.6]
  assign _T_1560 = ~_T_1559; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209918.6]
  assign _T_1561 = io_in_d_bits_size == _T_1547; // @[Monitor.scala 541:29:freechips.rocketchip.system.DefaultRV32Config.fir@209923.6]
  assign _T_1563 = _T_1561 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209925.6]
  assign _T_1564 = ~_T_1563; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209926.6]
  assign _T_1565 = io_in_d_bits_source == _T_1548; // @[Monitor.scala 542:29:freechips.rocketchip.system.DefaultRV32Config.fir@209931.6]
  assign _T_1567 = _T_1565 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209933.6]
  assign _T_1568 = ~_T_1567; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209934.6]
  assign _T_1569 = io_in_d_bits_sink == _T_1549; // @[Monitor.scala 543:29:freechips.rocketchip.system.DefaultRV32Config.fir@209939.6]
  assign _T_1571 = _T_1569 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209941.6]
  assign _T_1572 = ~_T_1571; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209942.6]
  assign _T_1573 = io_in_d_bits_denied == _T_1550; // @[Monitor.scala 544:29:freechips.rocketchip.system.DefaultRV32Config.fir@209947.6]
  assign _T_1575 = _T_1573 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209949.6]
  assign _T_1576 = ~_T_1575; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209950.6]
  assign _T_1578 = _T_1526 & _T_1537; // @[Monitor.scala 546:20:freechips.rocketchip.system.DefaultRV32Config.fir@209957.4]
  assign _T_1579 = io_in_b_ready & io_in_b_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@209966.4]
  assign _T_1590 = _T_1588 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@209977.4]
  assign _T_1591 = _T_1588 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@209978.4]
  assign _T_1604 = ~_T_1591; // @[Monitor.scala 409:22:freechips.rocketchip.system.DefaultRV32Config.fir@209994.4]
  assign _T_1605 = io_in_b_valid & _T_1604; // @[Monitor.scala 409:19:freechips.rocketchip.system.DefaultRV32Config.fir@209995.4]
  assign _T_1606 = io_in_b_bits_opcode == _T_1599; // @[Monitor.scala 410:32:freechips.rocketchip.system.DefaultRV32Config.fir@209997.6]
  assign _T_1608 = _T_1606 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209999.6]
  assign _T_1609 = ~_T_1608; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210000.6]
  assign _T_1610 = io_in_b_bits_param == _T_1600; // @[Monitor.scala 411:32:freechips.rocketchip.system.DefaultRV32Config.fir@210005.6]
  assign _T_1612 = _T_1610 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210007.6]
  assign _T_1613 = ~_T_1612; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210008.6]
  assign _T_1614 = io_in_b_bits_size == _T_1601; // @[Monitor.scala 412:32:freechips.rocketchip.system.DefaultRV32Config.fir@210013.6]
  assign _T_1616 = _T_1614 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210015.6]
  assign _T_1617 = ~_T_1616; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210016.6]
  assign _T_1618 = io_in_b_bits_source == _T_1602; // @[Monitor.scala 413:32:freechips.rocketchip.system.DefaultRV32Config.fir@210021.6]
  assign _T_1620 = _T_1618 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210023.6]
  assign _T_1621 = ~_T_1620; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210024.6]
  assign _T_1622 = io_in_b_bits_address == _T_1603; // @[Monitor.scala 414:32:freechips.rocketchip.system.DefaultRV32Config.fir@210029.6]
  assign _T_1624 = _T_1622 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210031.6]
  assign _T_1625 = ~_T_1624; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210032.6]
  assign _T_1627 = _T_1579 & _T_1591; // @[Monitor.scala 416:20:freechips.rocketchip.system.DefaultRV32Config.fir@210039.4]
  assign _T_1628 = io_in_c_ready & io_in_c_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@210047.4]
  assign _T_1638 = _T_1636 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@210057.4]
  assign _T_1639 = _T_1636 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@210058.4]
  assign _T_1652 = ~_T_1639; // @[Monitor.scala 514:22:freechips.rocketchip.system.DefaultRV32Config.fir@210074.4]
  assign _T_1653 = io_in_c_valid & _T_1652; // @[Monitor.scala 514:19:freechips.rocketchip.system.DefaultRV32Config.fir@210075.4]
  assign _T_1654 = io_in_c_bits_opcode == _T_1647; // @[Monitor.scala 515:32:freechips.rocketchip.system.DefaultRV32Config.fir@210077.6]
  assign _T_1656 = _T_1654 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210079.6]
  assign _T_1657 = ~_T_1656; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210080.6]
  assign _T_1658 = io_in_c_bits_param == _T_1648; // @[Monitor.scala 516:32:freechips.rocketchip.system.DefaultRV32Config.fir@210085.6]
  assign _T_1660 = _T_1658 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210087.6]
  assign _T_1661 = ~_T_1660; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210088.6]
  assign _T_1662 = io_in_c_bits_size == _T_1649; // @[Monitor.scala 517:32:freechips.rocketchip.system.DefaultRV32Config.fir@210093.6]
  assign _T_1664 = _T_1662 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210095.6]
  assign _T_1665 = ~_T_1664; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210096.6]
  assign _T_1666 = io_in_c_bits_source == _T_1650; // @[Monitor.scala 518:32:freechips.rocketchip.system.DefaultRV32Config.fir@210101.6]
  assign _T_1668 = _T_1666 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210103.6]
  assign _T_1669 = ~_T_1668; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210104.6]
  assign _T_1670 = io_in_c_bits_address == _T_1651; // @[Monitor.scala 519:32:freechips.rocketchip.system.DefaultRV32Config.fir@210109.6]
  assign _T_1672 = _T_1670 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210111.6]
  assign _T_1673 = ~_T_1672; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210112.6]
  assign _T_1675 = _T_1628 & _T_1639; // @[Monitor.scala 521:20:freechips.rocketchip.system.DefaultRV32Config.fir@210119.4]
  assign _T_1687 = _T_1685 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@210141.4]
  assign a_first = _T_1685 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@210142.4]
  assign _T_1705 = _T_1703 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@210163.4]
  assign d_first = _T_1703 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@210164.4]
  assign _GEN_75 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 629:69:freechips.rocketchip.system.DefaultRV32Config.fir@210183.4]
  assign _T_1713 = {{1'd0}, _GEN_75}; // @[Monitor.scala 629:69:freechips.rocketchip.system.DefaultRV32Config.fir@210183.4]
  assign _T_1714 = inflight_opcodes >> _T_1713; // @[Monitor.scala 629:44:freechips.rocketchip.system.DefaultRV32Config.fir@210184.4]
  assign _T_1718 = 16'h10 - 16'h1; // @[Monitor.scala 606:57:freechips.rocketchip.system.DefaultRV32Config.fir@210188.4]
  assign _GEN_76 = {{4'd0}, _T_1714}; // @[Monitor.scala 629:97:freechips.rocketchip.system.DefaultRV32Config.fir@210189.4]
  assign _T_1719 = _GEN_76 & _T_1718; // @[Monitor.scala 629:97:freechips.rocketchip.system.DefaultRV32Config.fir@210189.4]
  assign _T_1720 = {{1'd0}, _T_1719[15:1]}; // @[Monitor.scala 629:152:freechips.rocketchip.system.DefaultRV32Config.fir@210190.4]
  assign _T_1721 = {io_in_d_bits_source, 3'h0}; // @[Monitor.scala 633:65:freechips.rocketchip.system.DefaultRV32Config.fir@210194.4]
  assign _T_1722 = inflight_sizes >> _T_1721; // @[Monitor.scala 633:40:freechips.rocketchip.system.DefaultRV32Config.fir@210195.4]
  assign _T_1726 = 16'h100 - 16'h1; // @[Monitor.scala 606:57:freechips.rocketchip.system.DefaultRV32Config.fir@210199.4]
  assign _GEN_78 = {{8'd0}, _T_1726}; // @[Monitor.scala 633:91:freechips.rocketchip.system.DefaultRV32Config.fir@210200.4]
  assign _T_1727 = _T_1722 & _GEN_78; // @[Monitor.scala 633:91:freechips.rocketchip.system.DefaultRV32Config.fir@210200.4]
  assign _T_1728 = {{1'd0}, _T_1727[23:1]}; // @[Monitor.scala 633:144:freechips.rocketchip.system.DefaultRV32Config.fir@210201.4]
  assign _T_1732 = _T_1477 & a_first; // @[Monitor.scala 643:27:freechips.rocketchip.system.DefaultRV32Config.fir@210226.4]
  assign _T_1734 = 4'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@210229.6]
  assign _T_1735 = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 645:53:freechips.rocketchip.system.DefaultRV32Config.fir@210231.6]
  assign _T_1736 = _T_1735 | 4'h1; // @[Monitor.scala 645:61:freechips.rocketchip.system.DefaultRV32Config.fir@210232.6]
  assign _T_1737 = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 646:49:freechips.rocketchip.system.DefaultRV32Config.fir@210234.6]
  assign _T_1738 = _T_1737 | 5'h1; // @[Monitor.scala 646:57:freechips.rocketchip.system.DefaultRV32Config.fir@210235.6]
  assign _GEN_80 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 647:72:freechips.rocketchip.system.DefaultRV32Config.fir@210237.6]
  assign _T_1739 = {{1'd0}, _GEN_80}; // @[Monitor.scala 647:72:freechips.rocketchip.system.DefaultRV32Config.fir@210237.6]
  assign a_opcodes_set_interm = _T_1732 ? _T_1736 : 4'h0; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@210228.4]
  assign _GEN_81 = {{31'd0}, a_opcodes_set_interm}; // @[Monitor.scala 647:47:freechips.rocketchip.system.DefaultRV32Config.fir@210238.6]
  assign _T_1740 = _GEN_81 << _T_1739; // @[Monitor.scala 647:47:freechips.rocketchip.system.DefaultRV32Config.fir@210238.6]
  assign _T_1741 = {io_in_a_bits_source, 3'h0}; // @[Monitor.scala 648:68:freechips.rocketchip.system.DefaultRV32Config.fir@210240.6]
  assign a_sizes_set_interm = _T_1732 ? _T_1738 : 5'h0; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@210228.4]
  assign _GEN_82 = {{31'd0}, a_sizes_set_interm}; // @[Monitor.scala 648:43:freechips.rocketchip.system.DefaultRV32Config.fir@210241.6]
  assign _T_1742 = _GEN_82 << _T_1741; // @[Monitor.scala 648:43:freechips.rocketchip.system.DefaultRV32Config.fir@210241.6]
  assign _T_1743 = inflight >> io_in_a_bits_source; // @[Monitor.scala 649:26:freechips.rocketchip.system.DefaultRV32Config.fir@210243.6]
  assign _T_1745 = ~_T_1743[0]; // @[Monitor.scala 649:17:freechips.rocketchip.system.DefaultRV32Config.fir@210245.6]
  assign _T_1747 = _T_1745 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210247.6]
  assign _T_1748 = ~_T_1747; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210248.6]
  assign _GEN_27 = _T_1732 ? _T_1734 : 4'h0; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@210228.4]
  assign _GEN_30 = _T_1732 ? _T_1740 : 35'h0; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@210228.4]
  assign _GEN_31 = _T_1732 ? _T_1742 : 36'h0; // @[Monitor.scala 643:72:freechips.rocketchip.system.DefaultRV32Config.fir@210228.4]
  assign _T_1751 = _T_1526 & d_first; // @[Monitor.scala 660:27:freechips.rocketchip.system.DefaultRV32Config.fir@210262.4]
  assign _T_1753 = ~_T_708; // @[Monitor.scala 660:75:freechips.rocketchip.system.DefaultRV32Config.fir@210264.4]
  assign _T_1754 = _T_1751 & _T_1753; // @[Monitor.scala 660:72:freechips.rocketchip.system.DefaultRV32Config.fir@210265.4]
  assign _T_1755 = 4'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@210267.6]
  assign _GEN_84 = {{31'd0}, _T_1718}; // @[Monitor.scala 662:76:freechips.rocketchip.system.DefaultRV32Config.fir@210274.6]
  assign _T_1761 = _GEN_84 << _T_1713; // @[Monitor.scala 662:76:freechips.rocketchip.system.DefaultRV32Config.fir@210274.6]
  assign _GEN_85 = {{31'd0}, _T_1726}; // @[Monitor.scala 663:72:freechips.rocketchip.system.DefaultRV32Config.fir@210281.6]
  assign _T_1767 = _GEN_85 << _T_1721; // @[Monitor.scala 663:72:freechips.rocketchip.system.DefaultRV32Config.fir@210281.6]
  assign _GEN_32 = _T_1754 ? _T_1755 : 4'h0; // @[Monitor.scala 660:91:freechips.rocketchip.system.DefaultRV32Config.fir@210266.4]
  assign _GEN_33 = _T_1754 ? _T_1761 : 47'h0; // @[Monitor.scala 660:91:freechips.rocketchip.system.DefaultRV32Config.fir@210266.4]
  assign _GEN_34 = _T_1754 ? _T_1767 : 47'h0; // @[Monitor.scala 660:91:freechips.rocketchip.system.DefaultRV32Config.fir@210266.4]
  assign _T_1768 = io_in_d_valid & d_first; // @[Monitor.scala 665:26:freechips.rocketchip.system.DefaultRV32Config.fir@210284.4]
  assign _T_1771 = _T_1768 & _T_1753; // @[Monitor.scala 665:71:freechips.rocketchip.system.DefaultRV32Config.fir@210287.4]
  assign _T_1772 = inflight >> io_in_d_bits_source; // @[Monitor.scala 666:25:freechips.rocketchip.system.DefaultRV32Config.fir@210289.6]
  assign _T_1774 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 666:93:freechips.rocketchip.system.DefaultRV32Config.fir@210291.6]
  assign _T_1775 = io_in_a_valid & _T_1774; // @[Monitor.scala 666:68:freechips.rocketchip.system.DefaultRV32Config.fir@210292.6]
  assign _T_1776 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 666:142:freechips.rocketchip.system.DefaultRV32Config.fir@210293.6]
  assign _T_1777 = _T_1775 & _T_1776; // @[Monitor.scala 666:119:freechips.rocketchip.system.DefaultRV32Config.fir@210294.6]
  assign _T_1778 = _T_1777 & a_first; // @[Monitor.scala 666:166:freechips.rocketchip.system.DefaultRV32Config.fir@210295.6]
  assign _T_1779 = _T_1772[0] | _T_1778; // @[Monitor.scala 666:49:freechips.rocketchip.system.DefaultRV32Config.fir@210296.6]
  assign _T_1781 = _T_1779 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210298.6]
  assign _T_1782 = ~_T_1781; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210299.6]
  assign a_opcode_lookup = _T_1720[3:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@210181.4 :freechips.rocketchip.system.DefaultRV32Config.fir@210182.4 Monitor.scala 629:21:freechips.rocketchip.system.DefaultRV32Config.fir@210191.4]
  assign _GEN_37 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@210305.6]
  assign _GEN_38 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_37; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@210305.6]
  assign _GEN_39 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_38; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@210305.6]
  assign _GEN_40 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_39; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@210305.6]
  assign _GEN_41 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_40; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@210305.6]
  assign _GEN_42 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_41; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@210305.6]
  assign _T_1784 = io_in_d_bits_opcode == _GEN_42; // @[Monitor.scala 667:37:freechips.rocketchip.system.DefaultRV32Config.fir@210305.6]
  assign _GEN_49 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_40; // @[Monitor.scala 667:96:freechips.rocketchip.system.DefaultRV32Config.fir@210307.6]
  assign _GEN_50 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_49; // @[Monitor.scala 667:96:freechips.rocketchip.system.DefaultRV32Config.fir@210307.6]
  assign _T_1786 = io_in_d_bits_opcode == _GEN_50; // @[Monitor.scala 667:96:freechips.rocketchip.system.DefaultRV32Config.fir@210307.6]
  assign _T_1787 = _T_1784 | _T_1786; // @[Monitor.scala 667:71:freechips.rocketchip.system.DefaultRV32Config.fir@210308.6]
  assign _GEN_53 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@210309.6]
  assign _GEN_54 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_53; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@210309.6]
  assign _GEN_55 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_54; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@210309.6]
  assign _GEN_56 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_55; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@210309.6]
  assign _GEN_57 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_56; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@210309.6]
  assign _GEN_58 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_57; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@210309.6]
  assign _T_1788 = io_in_d_bits_opcode == _GEN_58; // @[Monitor.scala 668:60:freechips.rocketchip.system.DefaultRV32Config.fir@210309.6]
  assign _GEN_65 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_56; // @[Monitor.scala 668:124:freechips.rocketchip.system.DefaultRV32Config.fir@210310.6]
  assign _GEN_66 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_65; // @[Monitor.scala 668:124:freechips.rocketchip.system.DefaultRV32Config.fir@210310.6]
  assign _T_1789 = io_in_d_bits_opcode == _GEN_66; // @[Monitor.scala 668:124:freechips.rocketchip.system.DefaultRV32Config.fir@210310.6]
  assign _T_1790 = _T_1788 | _T_1789; // @[Monitor.scala 668:99:freechips.rocketchip.system.DefaultRV32Config.fir@210311.6]
  assign _T_1791 = io_in_a_valid & _T_1790; // @[Monitor.scala 668:34:freechips.rocketchip.system.DefaultRV32Config.fir@210312.6]
  assign _T_1792 = _T_1787 | _T_1791; // @[Monitor.scala 668:15:freechips.rocketchip.system.DefaultRV32Config.fir@210313.6]
  assign _T_1794 = _T_1792 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210315.6]
  assign _T_1795 = ~_T_1794; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210316.6]
  assign a_size_lookup = _T_1728[7:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@210192.4 :freechips.rocketchip.system.DefaultRV32Config.fir@210193.4 Monitor.scala 633:19:freechips.rocketchip.system.DefaultRV32Config.fir@210202.4]
  assign _GEN_86 = {{4'd0}, io_in_d_bits_size}; // @[Monitor.scala 670:34:freechips.rocketchip.system.DefaultRV32Config.fir@210321.6]
  assign _T_1796 = _GEN_86 == a_size_lookup; // @[Monitor.scala 670:34:freechips.rocketchip.system.DefaultRV32Config.fir@210321.6]
  assign _T_1798 = io_in_a_valid & _T_1776; // @[Monitor.scala 670:72:freechips.rocketchip.system.DefaultRV32Config.fir@210323.6]
  assign _T_1799 = _T_1796 | _T_1798; // @[Monitor.scala 670:53:freechips.rocketchip.system.DefaultRV32Config.fir@210324.6]
  assign _T_1801 = _T_1799 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210326.6]
  assign _T_1802 = ~_T_1801; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210327.6]
  assign _T_1804 = _T_1768 & a_first; // @[Monitor.scala 672:36:freechips.rocketchip.system.DefaultRV32Config.fir@210334.4]
  assign _T_1805 = _T_1804 & io_in_a_valid; // @[Monitor.scala 672:47:freechips.rocketchip.system.DefaultRV32Config.fir@210335.4]
  assign _T_1807 = _T_1805 & _T_1774; // @[Monitor.scala 672:65:freechips.rocketchip.system.DefaultRV32Config.fir@210337.4]
  assign _T_1809 = _T_1807 & _T_1753; // @[Monitor.scala 672:116:freechips.rocketchip.system.DefaultRV32Config.fir@210339.4]
  assign _T_1810 = ~io_in_d_ready; // @[Monitor.scala 673:15:freechips.rocketchip.system.DefaultRV32Config.fir@210341.6]
  assign _T_1811 = _T_1810 | io_in_a_ready; // @[Monitor.scala 673:32:freechips.rocketchip.system.DefaultRV32Config.fir@210342.6]
  assign _T_1813 = _T_1811 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210344.6]
  assign _T_1814 = ~_T_1813; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210345.6]
  assign a_set = _GEN_27[2:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@210175.4 :freechips.rocketchip.system.DefaultRV32Config.fir@210176.4 Monitor.scala 644:13:freechips.rocketchip.system.DefaultRV32Config.fir@210230.6]
  assign d_clr = _GEN_32[2:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@210254.4 :freechips.rocketchip.system.DefaultRV32Config.fir@210255.4 Monitor.scala 661:13:freechips.rocketchip.system.DefaultRV32Config.fir@210268.6]
  assign _T_1815 = a_set != d_clr; // @[Monitor.scala 677:20:freechips.rocketchip.system.DefaultRV32Config.fir@210351.4]
  assign _T_1816 = |a_set; // @[Monitor.scala 677:40:freechips.rocketchip.system.DefaultRV32Config.fir@210352.4]
  assign _T_1817 = ~_T_1816; // @[Monitor.scala 677:33:freechips.rocketchip.system.DefaultRV32Config.fir@210353.4]
  assign _T_1818 = _T_1815 | _T_1817; // @[Monitor.scala 677:30:freechips.rocketchip.system.DefaultRV32Config.fir@210354.4]
  assign _T_1820 = _T_1818 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210356.4]
  assign _T_1821 = ~_T_1820; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210357.4]
  assign _T_1822 = inflight | a_set; // @[Monitor.scala 680:27:freechips.rocketchip.system.DefaultRV32Config.fir@210362.4]
  assign _T_1823 = ~d_clr; // @[Monitor.scala 680:38:freechips.rocketchip.system.DefaultRV32Config.fir@210363.4]
  assign _T_1824 = _T_1822 & _T_1823; // @[Monitor.scala 680:36:freechips.rocketchip.system.DefaultRV32Config.fir@210364.4]
  assign a_opcodes_set = _GEN_30[11:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@210177.4 :freechips.rocketchip.system.DefaultRV32Config.fir@210178.4 Monitor.scala 647:21:freechips.rocketchip.system.DefaultRV32Config.fir@210239.6]
  assign _T_1825 = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 681:43:freechips.rocketchip.system.DefaultRV32Config.fir@210366.4]
  assign d_opcodes_clr = _GEN_33[11:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@210256.4 :freechips.rocketchip.system.DefaultRV32Config.fir@210257.4 Monitor.scala 662:21:freechips.rocketchip.system.DefaultRV32Config.fir@210275.6]
  assign _T_1826 = ~d_opcodes_clr; // @[Monitor.scala 681:62:freechips.rocketchip.system.DefaultRV32Config.fir@210367.4]
  assign _T_1827 = _T_1825 & _T_1826; // @[Monitor.scala 681:60:freechips.rocketchip.system.DefaultRV32Config.fir@210368.4]
  assign a_sizes_set = _GEN_31[23:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@210179.4 :freechips.rocketchip.system.DefaultRV32Config.fir@210180.4 Monitor.scala 648:19:freechips.rocketchip.system.DefaultRV32Config.fir@210242.6]
  assign _T_1828 = inflight_sizes | a_sizes_set; // @[Monitor.scala 682:39:freechips.rocketchip.system.DefaultRV32Config.fir@210370.4]
  assign d_sizes_clr = _GEN_34[23:0]; // @[:freechips.rocketchip.system.DefaultRV32Config.fir@210258.4 :freechips.rocketchip.system.DefaultRV32Config.fir@210259.4 Monitor.scala 663:19:freechips.rocketchip.system.DefaultRV32Config.fir@210282.6]
  assign _T_1829 = ~d_sizes_clr; // @[Monitor.scala 682:56:freechips.rocketchip.system.DefaultRV32Config.fir@210371.4]
  assign _T_1830 = _T_1828 & _T_1829; // @[Monitor.scala 682:54:freechips.rocketchip.system.DefaultRV32Config.fir@210372.4]
  assign _T_1832 = |inflight; // @[Monitor.scala 687:26:freechips.rocketchip.system.DefaultRV32Config.fir@210377.4]
  assign _T_1833 = ~_T_1832; // @[Monitor.scala 687:16:freechips.rocketchip.system.DefaultRV32Config.fir@210378.4]
  assign _T_1834 = plusarg_reader_out == 32'h0; // @[Monitor.scala 687:39:freechips.rocketchip.system.DefaultRV32Config.fir@210379.4]
  assign _T_1835 = _T_1833 | _T_1834; // @[Monitor.scala 687:30:freechips.rocketchip.system.DefaultRV32Config.fir@210380.4]
  assign _T_1836 = _T_1831 < plusarg_reader_out; // @[Monitor.scala 687:59:freechips.rocketchip.system.DefaultRV32Config.fir@210381.4]
  assign _T_1837 = _T_1835 | _T_1836; // @[Monitor.scala 687:47:freechips.rocketchip.system.DefaultRV32Config.fir@210382.4]
  assign _T_1839 = _T_1837 | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210384.4]
  assign _T_1840 = ~_T_1839; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210385.4]
  assign _T_1842 = _T_1831 + 32'h1; // @[Monitor.scala 689:26:freechips.rocketchip.system.DefaultRV32Config.fir@210391.4]
  assign _T_1845 = _T_1477 | _T_1526; // @[Monitor.scala 690:27:freechips.rocketchip.system.DefaultRV32Config.fir@210395.4]
  assign _T_1857 = _T_1855 - 10'h1; // @[Edges.scala 231:28:freechips.rocketchip.system.DefaultRV32Config.fir@210410.4]
  assign _T_1858 = _T_1855 == 10'h0; // @[Edges.scala 232:25:freechips.rocketchip.system.DefaultRV32Config.fir@210411.4]
  assign _T_1868 = _T_1526 & _T_1858; // @[Monitor.scala 700:27:freechips.rocketchip.system.DefaultRV32Config.fir@210425.4]
  assign _T_1871 = ~io_in_d_bits_opcode[1]; // @[Edges.scala 72:43:freechips.rocketchip.system.DefaultRV32Config.fir@210428.4]
  assign _T_1872 = io_in_d_bits_opcode[2] & _T_1871; // @[Edges.scala 72:40:freechips.rocketchip.system.DefaultRV32Config.fir@210429.4]
  assign _T_1873 = _T_1868 & _T_1872; // @[Monitor.scala 700:38:freechips.rocketchip.system.DefaultRV32Config.fir@210430.4]
  assign _T_1874 = 4'h1 << io_in_d_bits_sink; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@210432.6]
  assign _T_1875 = _T_1846 >> io_in_d_bits_sink; // @[Monitor.scala 702:23:freechips.rocketchip.system.DefaultRV32Config.fir@210434.6]
  assign _T_1877 = ~_T_1875[0]; // @[Monitor.scala 702:14:freechips.rocketchip.system.DefaultRV32Config.fir@210436.6]
  assign _T_1879 = _T_1877 | reset; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210438.6]
  assign _T_1880 = ~_T_1879; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210439.6]
  assign _GEN_69 = _T_1873 ? _T_1874 : 4'h0; // @[Monitor.scala 700:72:freechips.rocketchip.system.DefaultRV32Config.fir@210431.4]
  assign _T_1882 = io_in_e_ready & io_in_e_valid; // @[Decoupled.scala 40:37:freechips.rocketchip.system.DefaultRV32Config.fir@210447.4]
  assign _T_1885 = 4'h1 << io_in_e_bits_sink; // @[OneHot.scala 58:35:freechips.rocketchip.system.DefaultRV32Config.fir@210451.6]
  assign _T_1886 = _GEN_69 | _T_1846; // @[Monitor.scala 708:24:freechips.rocketchip.system.DefaultRV32Config.fir@210453.6]
  assign _T_1887 = _T_1886 >> io_in_e_bits_sink; // @[Monitor.scala 708:35:freechips.rocketchip.system.DefaultRV32Config.fir@210454.6]
  assign _T_1890 = _T_1887[0] | reset; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210457.6]
  assign _T_1891 = ~_T_1890; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210458.6]
  assign _GEN_70 = _T_1882 ? _T_1885 : 4'h0; // @[Monitor.scala 706:73:freechips.rocketchip.system.DefaultRV32Config.fir@210450.4]
  assign _T_1892 = _T_1846 | _GEN_69; // @[Monitor.scala 713:27:freechips.rocketchip.system.DefaultRV32Config.fir@210464.4]
  assign _T_1893 = ~_GEN_70; // @[Monitor.scala 713:38:freechips.rocketchip.system.DefaultRV32Config.fir@210465.4]
  assign _T_1894 = _T_1892 & _T_1893; // @[Monitor.scala 713:36:freechips.rocketchip.system.DefaultRV32Config.fir@210466.4]
  assign _GEN_87 = io_in_a_valid & _T_78; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207660.10]
  assign _GEN_103 = io_in_a_valid & _T_168; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207789.10]
  assign _GEN_121 = io_in_a_valid & _T_262; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207929.10]
  assign _GEN_133 = io_in_a_valid & _T_336; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208036.10]
  assign _GEN_143 = io_in_a_valid & _T_413; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208135.10]
  assign _GEN_153 = io_in_a_valid & _T_492; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208226.10]
  assign _GEN_163 = io_in_a_valid & _T_559; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208315.10]
  assign _GEN_173 = io_in_a_valid & _T_626; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208404.10]
  assign _GEN_185 = io_in_d_valid & _T_708; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208473.10]
  assign _GEN_195 = io_in_d_valid & _T_728; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208515.10]
  assign _GEN_205 = io_in_d_valid & _T_756; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208573.10]
  assign _GEN_215 = io_in_d_valid & _T_785; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208632.10]
  assign _GEN_221 = io_in_d_valid & _T_802; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208667.10]
  assign _GEN_227 = io_in_d_valid & _T_820; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208703.10]
  assign _GEN_233 = io_in_b_valid & _T_962; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208902.10]
  assign _GEN_247 = io_in_b_valid & _T_998; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208957.10]
  assign _GEN_261 = io_in_b_valid & _T_1023; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209012.10]
  assign _GEN_273 = io_in_b_valid & _T_1044; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209059.10]
  assign _GEN_285 = io_in_b_valid & _T_1067; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209108.10]
  assign _GEN_295 = io_in_b_valid & _T_1088; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209155.10]
  assign _GEN_305 = io_in_b_valid & _T_1109; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209202.10]
  assign _GEN_317 = io_in_c_valid & _T_1217; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209358.10]
  assign _GEN_327 = io_in_c_valid & _T_1239; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209406.10]
  assign _GEN_337 = io_in_c_valid & _T_1257; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209495.10]
  assign _GEN_349 = io_in_c_valid & _T_1342; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209615.10]
  assign _GEN_361 = io_in_c_valid & _T_1423; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209678.10]
  assign _GEN_369 = io_in_c_valid & _T_1441; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209718.10]
  assign _GEN_377 = io_in_c_valid & _T_1455; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209750.10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1486 = _RAND_0[9:0];
  _RAND_1 = {1{`RANDOM}};
  _T_1497 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  _T_1498 = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  _T_1499 = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  _T_1500 = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  _T_1501 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  _T_1534 = _RAND_6[9:0];
  _RAND_7 = {1{`RANDOM}};
  _T_1545 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  _T_1546 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  _T_1547 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  _T_1548 = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  _T_1549 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  _T_1550 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  _T_1588 = _RAND_13[9:0];
  _RAND_14 = {1{`RANDOM}};
  _T_1599 = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  _T_1600 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  _T_1601 = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  _T_1602 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  _T_1603 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  _T_1636 = _RAND_19[9:0];
  _RAND_20 = {1{`RANDOM}};
  _T_1647 = _RAND_20[2:0];
  _RAND_21 = {1{`RANDOM}};
  _T_1648 = _RAND_21[2:0];
  _RAND_22 = {1{`RANDOM}};
  _T_1649 = _RAND_22[3:0];
  _RAND_23 = {1{`RANDOM}};
  _T_1650 = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  _T_1651 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  inflight = _RAND_25[2:0];
  _RAND_26 = {1{`RANDOM}};
  inflight_opcodes = _RAND_26[11:0];
  _RAND_27 = {1{`RANDOM}};
  inflight_sizes = _RAND_27[23:0];
  _RAND_28 = {1{`RANDOM}};
  _T_1685 = _RAND_28[9:0];
  _RAND_29 = {1{`RANDOM}};
  _T_1703 = _RAND_29[9:0];
  _RAND_30 = {1{`RANDOM}};
  _T_1831 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  _T_1846 = _RAND_31[3:0];
  _RAND_32 = {1{`RANDOM}};
  _T_1855 = _RAND_32[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_1486 <= 10'h0;
    end else if (_T_1477) begin
      if (_T_1489) begin
        if (_T_1484) begin
          _T_1486 <= _T_13[11:2];
        end else begin
          _T_1486 <= 10'h0;
        end
      end else begin
        _T_1486 <= _T_1488;
      end
    end
    if (_T_1525) begin
      _T_1497 <= io_in_a_bits_opcode;
    end
    if (_T_1525) begin
      _T_1498 <= io_in_a_bits_param;
    end
    if (_T_1525) begin
      _T_1499 <= io_in_a_bits_size;
    end
    if (_T_1525) begin
      _T_1500 <= io_in_a_bits_source;
    end
    if (_T_1525) begin
      _T_1501 <= io_in_a_bits_address;
    end
    if (reset) begin
      _T_1534 <= 10'h0;
    end else if (_T_1526) begin
      if (_T_1537) begin
        if (io_in_d_bits_opcode[0]) begin
          _T_1534 <= _T_1530[11:2];
        end else begin
          _T_1534 <= 10'h0;
        end
      end else begin
        _T_1534 <= _T_1536;
      end
    end
    if (_T_1578) begin
      _T_1545 <= io_in_d_bits_opcode;
    end
    if (_T_1578) begin
      _T_1546 <= io_in_d_bits_param;
    end
    if (_T_1578) begin
      _T_1547 <= io_in_d_bits_size;
    end
    if (_T_1578) begin
      _T_1548 <= io_in_d_bits_source;
    end
    if (_T_1578) begin
      _T_1549 <= io_in_d_bits_sink;
    end
    if (_T_1578) begin
      _T_1550 <= io_in_d_bits_denied;
    end
    if (reset) begin
      _T_1588 <= 10'h0;
    end else if (_T_1579) begin
      if (_T_1591) begin
        _T_1588 <= 10'h0;
      end else begin
        _T_1588 <= _T_1590;
      end
    end
    if (_T_1627) begin
      _T_1599 <= io_in_b_bits_opcode;
    end
    if (_T_1627) begin
      _T_1600 <= io_in_b_bits_param;
    end
    if (_T_1627) begin
      _T_1601 <= io_in_b_bits_size;
    end
    if (_T_1627) begin
      _T_1602 <= io_in_b_bits_source;
    end
    if (_T_1627) begin
      _T_1603 <= io_in_b_bits_address;
    end
    if (reset) begin
      _T_1636 <= 10'h0;
    end else if (_T_1628) begin
      if (_T_1639) begin
        if (io_in_c_bits_opcode[0]) begin
          _T_1636 <= _T_1143[11:2];
        end else begin
          _T_1636 <= 10'h0;
        end
      end else begin
        _T_1636 <= _T_1638;
      end
    end
    if (_T_1675) begin
      _T_1647 <= io_in_c_bits_opcode;
    end
    if (_T_1675) begin
      _T_1648 <= io_in_c_bits_param;
    end
    if (_T_1675) begin
      _T_1649 <= io_in_c_bits_size;
    end
    if (_T_1675) begin
      _T_1650 <= io_in_c_bits_source;
    end
    if (_T_1675) begin
      _T_1651 <= io_in_c_bits_address;
    end
    if (reset) begin
      inflight <= 3'h0;
    end else begin
      inflight <= _T_1824;
    end
    if (reset) begin
      inflight_opcodes <= 12'h0;
    end else begin
      inflight_opcodes <= _T_1827;
    end
    if (reset) begin
      inflight_sizes <= 24'h0;
    end else begin
      inflight_sizes <= _T_1830;
    end
    if (reset) begin
      _T_1685 <= 10'h0;
    end else if (_T_1477) begin
      if (a_first) begin
        if (_T_1484) begin
          _T_1685 <= _T_13[11:2];
        end else begin
          _T_1685 <= 10'h0;
        end
      end else begin
        _T_1685 <= _T_1687;
      end
    end
    if (reset) begin
      _T_1703 <= 10'h0;
    end else if (_T_1526) begin
      if (d_first) begin
        if (io_in_d_bits_opcode[0]) begin
          _T_1703 <= _T_1530[11:2];
        end else begin
          _T_1703 <= 10'h0;
        end
      end else begin
        _T_1703 <= _T_1705;
      end
    end
    if (reset) begin
      _T_1831 <= 32'h0;
    end else if (_T_1845) begin
      _T_1831 <= 32'h0;
    end else begin
      _T_1831 <= _T_1842;
    end
    if (reset) begin
      _T_1846 <= 4'h0;
    end else begin
      _T_1846 <= _T_1894;
    end
    if (reset) begin
      _T_1855 <= 10'h0;
    end else if (_T_1526) begin
      if (_T_1858) begin
        if (io_in_d_bits_opcode[0]) begin
          _T_1855 <= _T_1530[11:2];
        end else begin
          _T_1855 <= 10'h0;
        end
      end else begin
        _T_1855 <= _T_1857;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_87 & _T_130) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock type unsupported by manager (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207660.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_87 & _T_130) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207661.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_87 & _T_144) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207683.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_87 & _T_144) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207684.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_87 & _T_147) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207690.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_87 & _T_147) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207691.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_87 & _T_151) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207698.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_87 & _T_151) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207699.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_87 & _T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207705.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_87 & _T_154) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207706.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_87 & _T_158) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207713.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_87 & _T_158) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207714.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_87 & _T_163) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207722.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_87 & _T_163) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207723.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_87 & _T_167) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207730.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_87 & _T_167) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207731.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_103 & _T_130) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm type unsupported by manager (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207789.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_103 & _T_130) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207790.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_103 & _T_144) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207812.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_103 & _T_144) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207813.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_103 & _T_147) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207819.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_103 & _T_147) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207820.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_103 & _T_151) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207827.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_103 & _T_151) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207828.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_103 & _T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207834.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_103 & _T_154) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207835.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_103 & _T_158) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207842.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_103 & _T_158) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207843.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_103 & _T_252) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207850.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_103 & _T_252) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207851.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_103 & _T_163) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207859.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_103 & _T_163) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207860.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_103 & _T_167) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207867.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_103 & _T_167) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207868.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_121 & _T_317) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Get type unsupported by manager (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207929.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_121 & _T_317) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207930.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_121 & _T_147) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207936.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_121 & _T_147) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207937.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_121 & _T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207943.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_121 & _T_154) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207944.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_121 & _T_327) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207951.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_121 & _T_327) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207952.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_121 & _T_331) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207959.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_121 & _T_331) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207960.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_121 & _T_167) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207967.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_121 & _T_167) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@207968.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_398) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutFull type unsupported by manager (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208036.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_398) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208037.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_147) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208043.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_147) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208044.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208050.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_154) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208051.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_327) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208058.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_327) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208059.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_133 & _T_331) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208066.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_133 & _T_331) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208067.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_143 & _T_398) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutPartial type unsupported by manager (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208135.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_143 & _T_398) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208136.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_143 & _T_147) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208142.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_143 & _T_147) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208143.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_143 & _T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208149.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_143 & _T_154) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208150.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_143 & _T_327) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208157.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_143 & _T_327) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208158.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_143 & _T_491) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208167.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_143 & _T_491) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208168.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & _T_544) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Arithmetic type unsupported by manager (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208226.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & _T_544) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208227.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & _T_147) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208233.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & _T_147) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208234.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & _T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208240.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & _T_154) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208241.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & _T_554) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208248.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & _T_554) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208249.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_153 & _T_331) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208256.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_153 & _T_331) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208257.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & _T_544) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Logical type unsupported by manager (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208315.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & _T_544) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208316.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & _T_147) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208322.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & _T_147) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208323.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & _T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208329.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & _T_154) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208330.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & _T_621) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid opcode param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208337.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & _T_621) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208338.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & _T_331) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208345.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_163 & _T_331) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208346.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_173 & _T_678) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Hint type unsupported by manager (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208404.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_173 & _T_678) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208405.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_173 & _T_147) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208411.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_173 & _T_147) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208412.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_173 & _T_154) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208418.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_173 & _T_154) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208419.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_173 & _T_688) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid opcode param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208426.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_173 & _T_688) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208427.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_173 & _T_331) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208434.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_173 & _T_331) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208435.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_173 & _T_167) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208442.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_173 & _T_167) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208443.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_700) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel has invalid opcode (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208453.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_700) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208454.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_185 & _T_711) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208473.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_185 & _T_711) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208474.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_185 & _T_715) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208481.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_185 & _T_715) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208482.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_185 & _T_719) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208489.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_185 & _T_719) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208490.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_185 & _T_723) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208497.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_185 & _T_723) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208498.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_185 & _T_727) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is denied (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208505.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_185 & _T_727) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208506.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & _T_711) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208515.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & _T_711) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208516.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & _T_715) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant smaller than a beat (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208530.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & _T_715) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208531.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & _T_742) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid cap param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208538.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & _T_742) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208539.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & _T_746) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries toN param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208546.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & _T_746) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208547.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_195 & _T_723) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208554.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_195 & _T_723) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208555.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & _T_711) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208573.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & _T_711) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208574.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & _T_715) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData smaller than a beat (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208588.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & _T_715) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208589.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & _T_742) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid cap param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208596.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & _T_742) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208597.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & _T_746) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries toN param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208604.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & _T_746) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208605.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_205 & _T_779) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208613.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_205 & _T_779) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208614.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_215 & _T_711) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208632.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_215 & _T_711) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208633.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_215 & _T_719) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208640.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_215 & _T_719) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208641.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_215 & _T_723) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208648.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_215 & _T_723) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208649.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_221 & _T_711) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208667.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_221 & _T_711) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208668.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_221 & _T_719) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208675.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_221 & _T_719) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208676.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_221 & _T_779) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208684.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_221 & _T_779) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208685.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_227 & _T_711) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208703.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_227 & _T_711) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208704.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_227 & _T_719) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208711.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_227 & _T_719) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208712.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_227 & _T_723) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208719.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_227 & _T_723) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@208720.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_b_valid & _T_840) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel has invalid opcode (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208739.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_b_valid & _T_840) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208740.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & _T_976) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Probe type unsupported by client (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208902.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & _T_976) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208903.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & _T_979) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208909.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & _T_979) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208910.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & _T_982) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries source that is not first source (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208916.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & _T_982) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208917.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & _T_985) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208923.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & _T_985) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208924.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & _T_989) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe carries invalid cap param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208931.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & _T_989) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208932.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & _T_993) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208939.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & _T_993) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208940.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_233 & _T_997) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Probe is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208947.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_233 & _T_997) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208948.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_247 & _T_1001) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Get type unsupported by client (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208957.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_247 & _T_1001) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208958.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_247 & _T_979) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208964.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_247 & _T_979) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208965.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_247 & _T_982) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries source that is not first source (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208971.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_247 & _T_982) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208972.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_247 & _T_985) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208978.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_247 & _T_985) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208979.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_247 & _T_1014) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208986.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_247 & _T_1014) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208987.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_247 & _T_993) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208994.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_247 & _T_993) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@208995.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_247 & _T_997) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Get is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209002.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_247 & _T_997) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209003.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_261 & _T_1001) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries PutFull type unsupported by client (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209012.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_261 & _T_1001) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209013.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_261 & _T_979) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209019.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_261 & _T_979) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209020.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_261 & _T_982) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries source that is not first source (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209026.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_261 & _T_982) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209027.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_261 & _T_985) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209033.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_261 & _T_985) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209034.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_261 & _T_1014) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209041.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_261 & _T_1014) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209042.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_261 & _T_993) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutFull contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209049.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_261 & _T_993) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209050.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_273 & _T_1001) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries PutPartial type unsupported by client (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209059.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_273 & _T_1001) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209060.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_273 & _T_979) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209066.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_273 & _T_979) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209067.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_273 & _T_982) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries source that is not first source (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209073.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_273 & _T_982) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209074.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_273 & _T_985) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209080.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_273 & _T_985) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209081.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_273 & _T_1014) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209088.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_273 & _T_1014) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209089.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_273 & _T_1066) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel PutPartial contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209098.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_273 & _T_1066) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209099.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_285 & _T_1001) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Arithmetic type unsupported by client (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209108.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_285 & _T_1001) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209109.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_285 & _T_979) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209115.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_285 & _T_979) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209116.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_285 & _T_982) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic carries source that is not first source (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209122.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_285 & _T_982) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209123.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_285 & _T_985) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209129.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_285 & _T_985) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209130.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_285 & _T_993) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Arithmetic contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209145.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_285 & _T_993) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209146.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_295 & _T_1001) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Logical type unsupported by client (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209155.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_295 & _T_1001) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209156.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_295 & _T_979) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209162.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_295 & _T_979) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209163.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_295 & _T_982) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical carries source that is not first source (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209169.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_295 & _T_982) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209170.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_295 & _T_985) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209176.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_295 & _T_985) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209177.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_295 & _T_993) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Logical contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209192.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_295 & _T_993) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209193.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_305 & _T_1001) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel carries Hint type unsupported by client (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209202.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_305 & _T_1001) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209203.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_305 & _T_979) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209209.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_305 & _T_979) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209210.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_305 & _T_982) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint carries source that is not first source (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209216.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_305 & _T_982) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209217.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_305 & _T_985) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209223.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_305 & _T_985) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209224.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_305 & _T_993) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint contains invalid mask (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209231.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_305 & _T_993) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209232.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_305 & _T_997) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel Hint is corrupt (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209239.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_305 & _T_997) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209240.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_317 & _T_1220) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209358.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_317 & _T_1220) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209359.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_317 & _T_1223) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209365.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_317 & _T_1223) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209366.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_317 & _T_1227) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209373.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_317 & _T_1227) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209374.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_317 & _T_1230) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209380.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_317 & _T_1230) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209381.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_317 & _T_1234) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209388.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_317 & _T_1234) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209389.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_327 & _T_1220) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209406.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_327 & _T_1220) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209407.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_327 & _T_1223) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209413.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_327 & _T_1223) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209414.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_327 & _T_1227) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209421.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_327 & _T_1227) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209422.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_327 & _T_1230) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209428.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_327 & _T_1230) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209429.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_327 & _T_1234) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209436.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_327 & _T_1234) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209437.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_337 & _T_1309) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release type unsupported by manager (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209495.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_337 & _T_1309) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209496.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_337 & _T_1323) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209518.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_337 & _T_1323) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209519.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_337 & _T_1223) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209525.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_337 & _T_1223) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209526.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_337 & _T_1227) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release smaller than a beat (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209533.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_337 & _T_1227) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209534.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_337 & _T_1230) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209540.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_337 & _T_1230) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209541.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_337 & _T_1337) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel Release carries invalid shrink param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209548.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_337 & _T_1337) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209549.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_349 & _T_1309) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209615.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_349 & _T_1309) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209616.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_349 & _T_1323) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209638.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_349 & _T_1323) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209639.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_349 & _T_1223) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209645.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_349 & _T_1223) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209646.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_349 & _T_1227) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209653.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_349 & _T_1227) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209654.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_349 & _T_1230) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209660.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_349 & _T_1230) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209661.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_349 & _T_1337) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel ReleaseData carries invalid shrink param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209668.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_349 & _T_1337) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209669.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_361 & _T_1220) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209678.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_361 & _T_1220) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209679.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_361 & _T_1223) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209685.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_361 & _T_1223) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209686.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_361 & _T_1230) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209692.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_361 & _T_1230) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209693.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_361 & _T_1436) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAck carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209700.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_361 & _T_1436) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209701.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_369 & _T_1220) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209718.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_369 & _T_1220) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209719.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_369 & _T_1223) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209725.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_369 & _T_1223) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209726.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_369 & _T_1230) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209732.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_369 & _T_1230) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209733.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_369 & _T_1436) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel AccessAckData carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209740.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_369 & _T_1436) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209741.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_377 & _T_1220) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries unmanaged address (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209750.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_377 & _T_1220) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209751.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_377 & _T_1223) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209757.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_377 & _T_1223) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209758.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_377 & _T_1230) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck address not aligned to size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209764.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_377 & _T_1230) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209765.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_377 & _T_1436) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel HintAck carries invalid param (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209772.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_377 & _T_1436) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209773.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1503 & _T_1507) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel opcode changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209831.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1503 & _T_1507) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209832.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1503 & _T_1511) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel param changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209839.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1503 & _T_1511) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209840.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1503 & _T_1515) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel size changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209847.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1503 & _T_1515) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209848.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1503 & _T_1519) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel source changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209855.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1503 & _T_1519) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209856.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1503 & _T_1523) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel address changed with multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209863.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1503 & _T_1523) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@209864.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1552 & _T_1556) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel opcode changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209912.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1552 & _T_1556) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209913.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1552 & _T_1560) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel param changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209920.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1552 & _T_1560) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209921.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1552 & _T_1564) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel size changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209928.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1552 & _T_1564) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209929.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1552 & _T_1568) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel source changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209936.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1552 & _T_1568) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209937.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1552 & _T_1572) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel sink changed with multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209944.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1552 & _T_1572) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209945.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1552 & _T_1576) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel denied changed with multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209952.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1552 & _T_1576) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@209953.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1605 & _T_1609) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel opcode changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210002.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1605 & _T_1609) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210003.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1605 & _T_1613) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel param changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210010.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1605 & _T_1613) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210011.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1605 & _T_1617) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel size changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210018.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1605 & _T_1617) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210019.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1605 & _T_1621) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel source changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210026.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1605 & _T_1621) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210027.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1605 & _T_1625) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel addresss changed with multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210034.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1605 & _T_1625) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210035.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1653 & _T_1657) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel opcode changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210082.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1653 & _T_1657) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210083.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1653 & _T_1661) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel param changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210090.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1653 & _T_1661) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210091.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1653 & _T_1665) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel size changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210098.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1653 & _T_1665) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210099.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1653 & _T_1669) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel source changed within multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210106.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1653 & _T_1669) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210107.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1653 & _T_1673) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel address changed with multibeat operation (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210114.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1653 & _T_1673) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210115.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1732 & _T_1748) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel re-used a source ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210250.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1732 & _T_1748) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210251.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1771 & _T_1782) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel acknowledged for nothing inflight (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210301.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1771 & _T_1782) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210302.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1771 & _T_1795) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel contains improper opcode response (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210318.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1771 & _T_1795) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210319.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1771 & _T_1802) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel contains improper response size (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210329.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1771 & _T_1802) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210330.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1809 & _T_1814) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210347.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1809 & _T_1814) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210348.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1821) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' and 'D' concurrent, despite minlatency 3 (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210359.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1821) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210360.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1840) begin
          $fwrite(32'h80000002,"Assertion failed: TileLink timeout expired (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210387.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1840) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210388.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1873 & _T_1880) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel re-used a sink ID (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:51 assert(cond, message)\n"); // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210441.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1873 & _T_1880) begin
          $fatal; // @[Monitor.scala 51:11:freechips.rocketchip.system.DefaultRV32Config.fir@210442.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1882 & _T_1891) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channel acknowledged for nothing inflight (connected at CrossingHelper.scala:30:80)\n    at Monitor.scala:44 assert(cond, message)\n"); // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210460.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1882 & _T_1891) begin
          $fatal; // @[Monitor.scala 44:11:freechips.rocketchip.system.DefaultRV32Config.fir@210461.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
